PK   mk�X1}��J=  b    cirkitFile.json�}]s�6��_��~ٍ5�"	޷nO;�;ݎ�lσ�C�϶�e鎤۶���� �$U�`Xw��1Ӗ�P��d"H$~�x����]�������Ǜ����2����~�~�O?�o���P����/�gO?�桯�����:��FH�dB�&3�ԙ��fà˼(�\��Z\����~w�AN��o��x��=]��J!T���h23�*�����u��A6����..�~\j�}QdE׷�ɭ��z�NhU֦�k�\�sq-�}���[F�5���w��{��b�]���Y}/}�̾v߹�:gs�"��́� �K6.���l\q]�9p�\����`J�B8�Ɂ�X��4±�L6�c�7�lǂo4���l�!��dC8|�Ɇp�$�v�!��dC8 ǚo;�v�!��dC8|�Ɇ���f����o;�b|�,��S�m�DW���&Ӻ�3#�<k����Do[U�]_!!p�_�r,�� Y�LÐ�Jԙcb�X��u�Ȳ�Fǆ��sK�<oF.w�q$ʾ��p�~���Y���Vwe#�N��;��+F��w��Z���(m��vn�ݏ�V�Y�6M��\�M�����B�;oFs�>gv~eF#vް:o�Oe甼j��o����1S:�D]+��v6��F���<J�{��{��{p����ٛ�w.���auŉ��rt ��0T�T��L��̌.DV��u���/r�K�������]���7�U�2Y�v��CQgu'�L��})�(��_[�N�,WG�>����j��b}a�ʂ���Ge��X_أ��B�/�QYp!���,���ڪ�zZ[����B�/�QY��ӵU9j�X_أ���εU9*��\[�����εU9*��\[�����εU9*��\[�����εU9*��d��-,�}�����[rb���������g��ǀ�J�:�=o����gLN�ȳ�9����;��'8�dw7�H��L�C;&����(oi����(dǤ�1B��횢�Q�j;�c��ON+vC;)�0g��1�w�'�+�k)��$���.(��������;�
o���T`p�1+��^b��Nbىk������Nbى�b+H�`��
63�H_&08H�������'��ƭ���Bt��B�JY7'�N۪�MQ�P��;al����9��с#8r���/l3HCɵخɅ�1E%4̒`~�o܎�/I0?	�7n������$�߸�4~�`~�oܼ�aa�I0�q�,?p���'���پD~ШB����P�Mpԣ�Q����4���.X~�oL/��w�޼�
(p���'��Ɣ������������X~�oL��`�I0�1,?p���'����5ئ&;��vS�:�R��AF�(pԃ�'���������������ٟ2��3	��$&���� �Q�jv(i�(��[_�LVF��$hC������M�Lg$;zN"��8VvԘ�z+;(;zba<BvPv��@�9u�쨱�<Vv�%Si���ِ��ݔ}��B�̴BhѺ��+�&��<V���z��2���ĝܠ����!�eG��V3�ʎQ+%`ee���C�ʎ��G.� ���_D�� X~�H
�o)�ni�"�	�쓫P�E�|~�E�s�"��ȥ7��GTX~Yz�!`���*,��,��W�T3���F$�������[T��T Z��ȹw��3`��W�ܻx��C,,����x���,,����x��C-�gOpx0W��a9��\�	� ��i|;� ��mX~i�;� �C�G�(r�<����_D��<����_D��<���{SX~i�;� ��2X~i�;� ��2X~Ki�8<�����_D��<�����:��ܳy)��ڼ�ϋ�F�|^�4���r��i{���+Ad$�y���LHXGF�f0�����ڑ=�p^��|��b��b�^3�.���w�+��{�+�)��=���
����~��+�U>�ӹ/�b=���i������������"�tj�P��K��yZg�O�q���Z��t͜�ux�'���m^�HT$������<c��S�B���1)(2!�1�+����+��LR��8� HR�H;�Ĥc�}GHv�x�Y���v�X���X��g�g�PˋZ�j�2z�4L����61�2�Ã����HL��X���Ɇb�L.��6CV
SdF��ݖ�9H��e��i�!x�2�h~h�!=9t�1��y��Ċ<��7�3	y	D,�(}ƓC�6�~�y�w�����t#d��/c�B���q�R�?�8�~^p$�<��H�yx�����Cp���!8�b��+(����/�����ArC�)?���2�s�h����)0��u$�̝f7�xse�2"īa���!]�����E�1�'M�tLwy6 �NT������������æ5��߉�S�rO@�Ze�j� MkEFG ;T-��B1����L�c�Q�& ����x��H��:�H�.<�H�Q�H���H���HL��D���b�8�����8�����8���ȁ8�����o����@�`\�L8
IL�i N0+.af�$�,:�c	��
f�QHbʸq��q��($1e�8�츂�q��2�@�`v\��8
ILY N0;�`v��D<A�m|��#Po�Z�m�^�ܴ>��B�m^������1�6��T�B��h��ئQ�tZg"2�6��|�	H���m\j�%���6�DF  �
yKd�{��L��J�59�B����h&'��!��P���0N0ӍB"���wga�`��DZC!�h�q��pi�\J�	f�QH�5r�*'�G!��P���`�`v�DZC!���q��qi�\��	f�QH�5r'�!�ӎ�_BQ��)�����տ�!��1�\���@����_����H!F_�
1�Q�r�/���5W�0��E�@����������!hRp���H`^c_�1��sE��犐�8"��)���a$0/�G�5W�f0���1v`^R��_�������b���iB�$l.�(�wH�®4q�w3Ѧ	��B��&��n�	!M����µaxX�lӄ`I�.���E�6M�����_xX�lӄbI�.\
��E�6M8���axX�lӄdI�.\&��E�6MX�����`xX��B��,	ۅ���H٦�˒�]�U��m�-�4q�w�)�4qY����a��M�%a�pS)�4qY����a��M�%a�p�)�4qY����g�H�~��"�4q�w���i�X��3�qd�Qa\��W_�}��m�a�3I���B�kd.%5�7�\#�jq�����S�I��P&'�k
�����@�����H=��D��1M��<@��\�52��G�52�2����L<*P�)�F�'Rk$�kdC-;�D�)�.�'�Q�rM�5:?�\�!M`�&�J�6>?�\g"�lE])�.�'B��4�Wl����P!m��+6�o,R�i¯$l��w�"e�&[`�	i��،��Wr�lB
����;`��M�6>?�\'�l�DcI���'�����m��,	���Dr��4�M�%a����WH��f��k:��ZH��f��E�6M\��m|~�X�lm����b3�v�"e�&.K�6>?q,R�i�$l��w�"e�f{,	�����H٦�˒���O���m��,	���D4,R�i�$l��w�"e�&.#�}�b4V
����E��AUY��_�������MJ��l$J�:l$J��k$J�k$J�;G���F���˱�(�J��(�ڟ��b����}.R?�` �p'�w'@,F�C��ca0*���Q�P%�X���'&p�N,L���X���6�0��hbaw���6�+�ca&-��r��9j����X�I��۷cg]�-֛�X��Sf��Cf�ͪ�0Y#T��N��W�6�P�֌i���ِ�E�MV�ƙi�ދ��t}�ͅ��ɥ,��U��}�eƶ}�(�g���j#����Q���DBQ[�6	EozXMgU�LV�]�Ԯ���ͭ�t�v��T��cDB�#ʶAA��"Jm��/�����ʬ��>�Vemʼ�A_((r�l�PԖ�$��-�IB1[6����\V�m���Ȍ*ݘK錖-d�ka�r8�Q�ho(�1*M��Q�� ��T��T%��E�v�Qg뼑eC�u$���$A1[cDB��ʦ+NB���I(��8	e��iݦC���`h0
�*a��M��(4�|+*p(EQ�ʹA����s�V�Y�6M��\�M�fQH(rK�$�M+3T�T���I��ֺY]�u�k�����G���f�H(�=j�)���ܔ^;�����T���U�ڣ���P6{DB9�ѯ������S��_���6�J᱗w�������_��� ��
a:��F ��oa:\�a:\�a:\�a:\�a:\�a:\�a:^ߋ1�8��3�0�-a��t���	f�%�x�����b8�췄p���^'��0#�B:^ߋ���
f�QH��{1�p�7���q��(����N0;�`v�t���	f�̎�����b8�츂�q�����B=��b���PSQ���.�&�ѶѥV�B1�6��:T(F��Z�	�h��Rk�m[j� #������k��L$�j��6�nV>�uQ`�`��DZC!��q��oi�\��	f�QH�5r�'�G!��P���a�`v�DZC!���q��qi�|n�	f�QH�5�9Q'�G!��P��a�`v<�ςW��z8n@]�b �
�p� (�\��H��Q�F�5ׅ+ �ꓠQ�rM�u����$hT�\Sp]�b "�.	(�\��H��I�F�5ׅ+ �ꑠQ�rM�u���Z$hT�\Sp]�b "�	(�\��x�i.�h?ƇOr%a�t� )�DaW���/��E�6M蕄��pX�lӄ_I�.]1 �E�6M����pX�lӄaI�.]1 �E�6M(����pX�lӄcI�.]1 �E�6MH����pX�lӄeI�.]1 �E�,��˒�]�b ��m��,	ۥ+�H�&�K��E��H٦�˒�]�b ��m��,	ۥ+�H٦�˒�]�b ��m��,	ۥ+�H٦�˒�]�b ��m��,	ۥ+�H٦��b�R�xƑ�G�q��O�G�52ȉG�5���Dj�o�F�7�,�$rM�5:?1(�\���g���52���N"�\���Q�rM�5:?�z=�\#��Q�$rM�5:?1(�\���5��52���H"�\���Q�rM�5:?�\�!M`�&�J�6>?�\g"�lE]�®4qWl��X�lӄ^I���'�E�6M���m|~�X�lӄ`I���'�E�6M��m|~�X�lӄbI���'�E�6M8��m|~�X�lӄdI���'�E�6MX��m|~�X��B��,	�����H٦�˒���O���m�-�4qYl��X�l��eI���'�E�6M\��m|~�X�l��eI���'�E�6M\��m|~�X�l��eI���'�E�6M\��m|~�X�l��e$�'W�+�PM�ڢ�̠��V���uc�tc�&%Pk6%P6%P�5%P�5%P35%P�4%P�4%PI4%P�3V�@ʋ��P��X���J���`48Tp=�á��0-���`���j��`�8T�:�š
ѱ0-�a��u1Z�7�X��Sf��Cf�ͪ�0Y#T��N��m������*��]/�!��웬Bd�B���t}�ͅ��ɥ,��U��}�eƶ}�(�g���j#��ns!�`�lʶ�i:�:e���J�vE�՝h3�]��T�^���m�)(����)�R�~�"+:��&�2���:�UY�2�mC�
ʶ�PP��������DBٜ�L.��6CV
SdF�n̥tF��̵0m9l�	es��� ��T��T%��E�v�Qg뼑eC�u$�M}!�l�	eS_H(��BB�tbH(�>	eӅ!�lz04�)/F{��IF��I̦;��(m�� ����9�U���h���M�ʦض2$��q"�l�P	SI�3�;w��Bdu!T6ԕ��.r����P6{DB��QSwM�7}6n��`���i*s]و�S-�s �l���rڣ_/ݟ?=]�����7�O������x[��׾���������~����u�Y�;���VM��RU����}]���Y}���肵dx4�8k=~�s�a�Ø�K�gL�h�] $3��I����d2�q��92Q���{�g=]�.yOW��+��5���t�{zp򠮕��γ�)y�Sz�T;9��=�T�v�8��x}�A����=�Vy@.�\���+ɤbH�qq|��΋.8TB����ԕ���K �"=��$I��£�V��g����0n�4����볲�%�~�6�{uۦ1E��}��v��Paڎy
,��
M��[`yO���3����t��_𞮃�"y�_E������K�������6�y�m���i��0a�d͋�Hr6�E������a4��7~e�|Hھ=/ޠ���5w�7�S*��$Ĭ�4s(1�%�4F��	�1���]V�9�y�H�u��e�(�g8y@�'BJ�.1'̀��&80�x	�y�scX�S=�[@[t���;��/Γ��&~bzϛ���st`T k~W����1����U7b��m��zvy@��[1�x�+i@��V,&k͞�N���⚵�.���oY��&�	qi~�o�d�u�-�iz�[�2���1/���Ǽ��[��0,ek���&�y�}��Q���p�w���w�Rv�o�b���tf��� �5/���L��
��¿?�$l>!p.���+%�T q-��ۦ��%����.�_�77~�=Z�ة�o9d�A� ��$ ��@ ��\ ��x ��� �� �����t�B�X�W������1�Om��q����MN9��;�2z�3|F�a�m�l���޵���ۿk��}����s��}�2]3O�@80���̛�G�3BKx���) �C* ��* �#+���osry�y�y�%�i����}��^$\�@p�"\S���4����'�V�߂BB�jo>d�17ׇ�WK��G<��QJyz�m_.Oo|���b���}\]8}�>���ЇS*Գ�)��Ŕ���b�@�z`qUC�s� �<����r[��m�P(��R(�NT�	0VB�;��J	�1K�P�O[��]��ܷ���s�Ӡ`��?�'�>���M����O�BL���T���(���(d���HW���I���gJ1�d��� ���t�ٚ�.l��oq�5츼	����Y���l~̒)"�ZBD�#˟���-0�q��爲���x��E�Yﰈ�&zX���6�M�ſy�坎g.W�W@��V@?���y)��_)޲H�ۡ�����E�G��n�����������q�O�ןn������A9\�{�MK}!��	�����|R�'
ب�OJ��B'ߨ>���I�R�>)6���ze�`C��X&6����e�`C��Z&6����e�`C��U�\����v�<��pY/�Cn���`c��u�\ +*f��!�J?| K*����x �)�� �S>ƘYp� �T�)C��>�< �T�)C�%?�< �T�)C����< �T�)c�� � �S�����Y\��u���.@޽�H�Jଯ��S<R��5�IN�H�*���Ϲ{�B�x���l)� �G*t��HjͰR���6`ͬY�!�WȉE����p��^�ְ�.m�)��y�B��f�����@� �0�|��%��&���16��< fwuy��O���|��%����� ��ccl,1Py ���� ����.Py ���� ����.Py ���� ����.�� < ������@N��c�5��N�&�/EË X��^�j�4��l�J(?�ć7Z��f��[�]f�Ն�0x ]����Aĩ�ک7���uKW�t��7`q�uq*�i�`�ҧ��~g~����� ����R��F/փg�b/ɞ-]�.S�%X;K�vb�I0?qm��`�a�I0?�(���1O�Uo7����3�����������`��п%�����弲9_����K�C�sn@��|�\	����ae~��q��𮻀bd�v��w
��!:�3��2�F�P���3��#0C��;����F��0C�f(��cbd��$����\��b:�3�h��>?Z���P��9
h�wj�[5�8E����S�%����!:N3�h����`d��S�%�ᘓ��!:N3�h��+2������p�{f��y�h�U�M.��J��k*A1Z��b������ �r�����;$Xu�"2��� ���D�0�����'rX��.�_D��%X~䈂z<,?,����x<����"rШ�R��#G��c!�����!���BJS��b_eW��̻رt#r��� ����A�jˏ=POL��巐��Ã��/"ˌ|T�|�c0Ø,3�v����RZ�l�
�^���E�[|�3	�r�w�c���s�ȵ�Z��e�9\; 12D�3>��*���t� Ĉ�c8� �%��A��)�aL��Z����0&�\7-Cttf��F�y��!:�3\�A�yV��z��@̒8:�3�II���!:�3�II���!|o���v bd�j�cR�v bd�j�cR�v bd�ާ3�II���!:l3�II���!:l3\JIbd�[�c��v bd�[6�^Ǘ+�PM�ڢ�̠��V���uc�tc���^Y���{�#�Q���W�0��������ꃑ�/7r�"�����KNK��t, W]�B�����P��r����5�ર_I8���~��X��uE,��%�x[�?��m]���u�B,�օ	�x���X��m����ř��o�ǎk��+v\��Sf��Cf�ͪ�0Y#T��N�酫bd@aIp��)��n��l��;�׳�^�ʲ�zQ�Y�7]fl�g��y&�Z��0������D�[�m��0$8߲ɐ%j:�:e���J��E�՝h3�F��K�D!�dr(p#�(p���۔��C_Yѹ���Vfu=���᪬M�׶Y��9�Β�.l�����#�|م,8	ΟPC��ϧ*`�L.��6CV
SdF�Ne�t���̵0m9,�l@�Hp#�;ҍ�>;�	���;P��w,���,	��;�P��*�߯D*�߯*�߯�)4U\��h +~`�l�Wނ�x4��H$`�ix�H`spEQ��yuֹ'�s��V�Y�6M��\�M�t�a���|ۤ�%�-ئ�;T�T��L���6�Y]�u�k����r�y
��$���������P4uה}�g����6Ϝ#�2Օ��:�.y;�������{A�[�lq����+�Mw�t��/��rA��.�{1��8ߌZ7vw��8(�M��3�8�L?%�L���L!��M.��L���bO���CM~���MN��DNFg��d<MR���f��F�� ��%.;�%��~H��Hq��C� (��Y)��qu�8�#ʫ��Hw���NdN܏
5��n�*������kIy�<�Ry�������!��<swEY��.FN߹���ᵻ�Ʒ���Й��P�/�މON�ȍ�m����:#��b֚2ˍ�{���a�(~L���fgX˭i�39�3�������ߛ����D��ĥD�3%�3�m��rm����Z �fnHKiK�~o*foX��!�A[v�:#�3�M� �1�ߗs�����-��f�]�aǪ���٩ ;�>+�(�"W�wVX��'�}v%�St�S�;|���7r&��N�J�;#��a���=��yD�|jU8NgB[��-(�3A'�zq �3��W����F��M�+��[�H�!�57�P�$Gܱ����dB�"�(q�=2Zp�0��y:4gc�������w�j�{r(���,vb�\ȟ$�I���;�Cqџ7�[�9l�9�eAC:G̗`�3[�B:G̫a���6���<�jN8�� �-��jĭW���#:$:�N.�]��5���v����LԜ��"��?�����EN6������o릿��Ĭ�/��?�_��W����Rǯ���>~�����+��������W��Uy�����ǯ��Uu����]�~��3{�ӗ����_>�J��}�~��s��;��S�<��*H�˸�\���)��4�/N�,N��S=�N��SϿS���s���?��?��O?����H?����H?����A?��^���)�y��yjA'�e-}Y��1��闗���z��������>� �D�����d���n����y|�6ǻ��Z�?�sV��]V����*[�e��u������k)����>�yF5m�\ ���W���tn��H�`����o� ��s��at2*�����lmUTn��eu�[Y��L���YG���~xS\L�r7�*��f����91"�E�M����a,�����og\Z��U�<��qf���\_�q��m����q�])UdҌn�� �Pd�)D�������l���Zd�P���M���j��\����<��B�n���o܄YU}����=Ÿ��c+����,��FYW�r�F���U(Y���*������heQ��U�<��|�&͝Z���*�.���#i�|E��9��-x>n/N���O�c����������~J�������їpo�������_��?��=~{y������_��^��h|��qݼp=~���p��qݗ���_no���峇��>�<�UO���?�w���}���?�8mv���tsw`�8��������[��+�_���ʝGR_��JwMn���ȉ�4�u��j2۸��˼4f��/�K��8!�ˋ��ǧ��= ���./�nJ}`uqx�o���8��:p�_#���V������������sg^�V'��ϋ���I����\�~�b�׿��窴�o���ߕ~�[��ϵ:�\�|��|^�|nO>�^?7���C_�������s{�y����_ǿ���������FE�su9��v���/&��p�����������.n��UؼS���Z��v��L]�ɼ�r�v�+��}����{�����ۯ�m��)��Mi��Rg��tV���tۗN�ߎ�?��iL=*T6�ةo�f���fZ�zt���/����㧧�ת�]��N��.��#�W�êE�7������ǯ���!�������ړ/����N���$��L��ɣnn�l�5�{7�ÊFg���~x�������k������u�H�q=A�u�J��J۔������)7��޺����ɧ��t/h[�茪ձ���c}���`;�g���a� ����� �Ç��?��tw?���៞�������~�u����_/�q�h�������}T��u��%�l�����錛w���ZV!��!��(2�t����s���uf��r�K
V�]5Zeλps�q>F%s7�Ճh��=�A����{Zۏ)�}1�L�LT�MtVw.:_W���.�~ӽ{�>}����/>ܽ{�/���=�����߼[����/�=ݿ{�t���Y������_���n��q~�o�`��}��w�?�������Ӥ2�_/����z��1��ڛ{�h7Gk����o�>u7�/�Ʌ��W�)w"�z
��|w��ç��w_�u������t����qz9����s��+#�����=��ˮ�U�;��;M�sgR�R�΋/e��}iʖ4Փ��S}w��7��D���<LQnN:~%���;O���.%W�o��'7{�E�h�7뇿}���>nԯ�_H�_��1Ua��k(k]7gn/�N����L�<���t�⦞�/��$}���r��R奋#]��l�t�:�ϕ�?�����=�o]�"F����w�}�]�s�����d��䩯��T\湹�,��"����1F=W;�O���,K=z��4}�GM΅c��r���ꠧ�8��,��N<��:p&��v��UV��t���N�q?�M��k=Т6�	B�VLQ[&Ks��aFK~�.��ߙ��N�R���-�i��⭔.
�%-�L9��h�S��]זj�n��&SE���F�0��eSԝ�ME�(g�*7.q:�c0.e^^�\�z��8]N�����Ӆ(�y���,�2��'���\Ϭ(���Y)�a���J���xx��g���M����lh:]���\��B=�u���]�Z���jѐԍtR��|�\��IY���ȯr�F�h�e	��VVWFm+��B]9Eֺ8Z@m�V���Yg]t���r���2Q��霫V�K5��$QR�b�̫�z��U����eU�ǥ�2?�r�˼����5'_�N2�	�<~Y�|'��\ZS��y��;�_��JW��4�;A[m�|�&���E���N-��Zh��j���3�9kQ��C[�=eC8��u^c%���ίwO�gl�f����\�7S��	�M��f�v���DU��x!*7x��r�G]�	7�y�>=�x�/E%�Vn�)�΅�RY]�<+{��ޚ������� /a��Fkq�2�Q���2���`��k��k�r��ׁ�������՟���|�_���\��͟��l��&��̌�G�|��O�O���E���no>~�<�_ߴ�y����/�>.U]4u���>��뾸��?�5_��ۼ��w���z�_��u{��<�zy�\�3Z��_�=a}P�u�����77��/��|��Ql��N�}q�ɽ@�����Fo6I
���*�jt"��\Hi�)�Ԧ��R��&�V�mԸ�Pe�l̸���BumtY(A�HG�mB��C��S�[^�.�q)ǔW���*�O���E.���r]��Q��1�.�ͥjd[Hّ��T���.�i��MS2�����;N�/_�s`��8�����H9�1�PΙ�tcye��)M�!U㠩�r��v���9��G��y���I�<H�9��j\�]l0���_�f�����_|�O��.�[���+-)�r����������U�́����2;|�b��czC���_dZ��W1�i�۵V� �}��M������ꕔfJ�������SKr\���WL����s��DW�~�wxI-���z��/7������q�/�e��vZ6m�N���0Ӗ��փ{���R�(n=�	����$U���tl?��8�V?}?a���Ç�1�������L&�q������NV/��9�V��K���V����VcԿЪ���Z}�뇋_�N��ח_N�իL�^�J�իL�^�lc�K��k��.�Dq�1��\V¹zy����Em-W�kG!���뵥R����OM�>�+�Xׯ}\#j6pί'�$��*gF��j�є�وj��P���R*��*]W�����b+)���Gl&�ZR)��=�^W��f�k�͖5tz�Q�5T͢L��m�.=�ACfq�*`�̎VfQ����FT���JG+,�R��V1�*S�Fq�J.*�gi�r�l;����͞����	��+�Z;�N��ک]�������Aq�[���]u�ߑ����S:Z�ٔ:G�vT�*�v筤^���S���32f-��(h�t:M�h�w�JA��
���I6�U��Oә��FT��JG,%�R��!j�P��}:o%e�1*�4;M���F!߾�e�'4b	�<ڈ�[�$˒̓"�������f+ŤF��͔�VA>�ΑmXU��Lج�YTL�νzR+��>q~����\ڪҍu���~�{��.�̙�-ݾ��"�k�]�;Z�l�,���"��o�v�&Rj���[��(�U;Z��ͧ�#��V/go7ԩ��h�Z,pcT&�:%zgT�
;mI��f��X�D?�P�V�,�T~6_�[�6��T�Hw�$�;�%���T���:o���%��B�B��tVvMV�
h~�����r�mN�f�BvE�l�y+��G��O��VD��jG�*��amD��缕{.E�����u�l`q��J�lz�]J`H~�!�C�O�ԇb92;_� �"[�7S:��m)��ly"�2�.`yf�ybҚ�^� %�v�ފ��/��R�]\)9����sZpH���c�W�@lF4!Q'1h�b�B�<���tc�b�J�=��f�̀��]	I�]7D��;�*�l����.ηO����Q��V˩G�EGR#�r�rѮ�*��O�vEpj��X��xY��!����Z�ryY؞O1�VI�l��[Ū���DpE���X�y��)^U�t�r�U�<V%�'+R+�y�Vٶ�a�2\�����J�ڬ��>��>��e�2�g���4��=��v���vrJ]٘�vQ�J(-��8 �Z�1�����ءj���<�d�)�D�O[fǐB��Y�d�jO+r2ś)�^򔺂5,�� =U	C٣:-,ьhX��y�zI<а��E�K�O[
��RP|���=�Ѱ������=��d]��]�����$��8)aӌhX��o��+�s?E:e�h�R�Ӗ�汔$_��ӊ���f�Bz[���ukXv�z�2,�f˙'��c�K\I%J�q��|~gI%:U��{q��S	�?��Ak*�4;QC\��+�F����bot�iTg��\uHeB���sOijMT
ډI��C�7b{��E�0�D���k�����|v(Ծfg�e�����׽v��n����#x��Lk�E��2�<�x�r�|@Q�j��e��S�`R!�6oEٝ�JW`��]�
-{�3� 5�S[����0lՉ��<h�Ք]�(F^WZز��^/�1�vsk�D9$����HP�����Tcߚ�|����R���l܉͞���5���gãb`��`�&R��,t�6�)��b�m���rֱ곷(uU����R�^��f�@	�Y�@=�y��Y�4m҈���wz�T�Y�|g��:�|UyΛ���{��fD�7��J��'���'�*r��[���K�.ڊ�����͒X҈`-��iy"��g��4��}O��3kFۆ$6Kj�6ڈ�����=@�
T������U��8z��K���NTg��*ɜE��^�Rs��{lc5G���h�>�D����P'�N���N��cR�D���tF��P�ԉ�������S���3�/�=k���5�� 5J��@�'Ng��DpE&%�]���C'\g������Y�$�ICA�����47\�j�@7VmH�+�Te�w&gm�XZF	v�H�Y-�K0t��o��*�Ѫ��4u~���rU}��V��o���U��%я[�&����O�������T����|��Ԭh�y�'�UhCl����E־гi�M�q1?�;r�,�w��I��wf�BN�x����퟇�����������J����w��[}������_=�?<�l������PK   �h�XWC��)�  � /   images/093f54e3-331f-4155-80d0-fca9fbcaa25c.png��	8���?>ҡ�)�T�9�TBC�,5��A�(Kd��/�q��2r�fP1ɞ�0�Q�
���=�k�}��~�z���������{����y��{�_���ǣkښ<?���\�����.��~r��>9��"�؉���]���u���K7�0ؑw�v7����0�='k��-�;0��v��h�[�wN;��ď�?��
����O�h�O� ݯ{~bz9a�.n���(��@�n�OoF�������_��v,ȋp�qW,��!��U�Է��N_�W��+��ޫ�}���.}�s�����}2lTSr��i�� C�s���sJJ��i%������鮋��?�������� T�źȜǾ�'w��A�t�+��OhEz8Ϥ�/e�>���e�%���%O��'�3W�L�����TV^&�o^����{��b0���.+Ű	�~�8�O�m���z�K��n��矌�t��d�D��`���JJJ�a��8�]\o7��N���;�Y��Kxrt�
Q����G��jm$M�KBS�='{�VVX+���i6=�˯�hT��_�1g���a��p�ݥ���6zC�*��4?,V����U�\p�{�3xc�w
C���\�"��	Z6�{��O$�O�(����Wj%�X����K���}�u�=���'�5�^%U_��~��!a�@G����1���̦a�w��W���4�8�$,䄞/���v�G�����^�-^CY�	�S�	�n���!T�17�!~,){$'L#Y'I�c�*1��9H	���|$��~��P�M�P�?%ͬLZ����{�OY�'L�oUۿH�H��������e%���OƯ���CkBW���Ou����Ƥ�n=`���C�\������Ŕ����ORŖ� ���۟��(����򣂒WP0;��e�*m>���G]�
�i�jl喨4eX���[\Hk��������6��ņ�\�B�m;�=��U�C�89ݻW���sv�~7%�f�J������n�2�oQ����u���^ۗ��% �5��£9�Z��;��� �1����p�`�g��7�Zt��nf��J/���DvE�.�5�b�`=ۥ��"֛�����K��ͫ��C��zCq'�sN�z�N�����j&ӟ�Fs�/��!�;�p�ԓ��8�L�aOǆ�{�����BT�}��dPTbߘ{1�K� ]���`��8�6JqSV�K�O���0�`u'��oB-¼�E��a��+��G���s�.��/�2��|cB��6]�`�2{��TW��wAR>ڦ�ªIϕ�s��}�z+/��Ra@�;�b�.NӍ�;n�`y�O�X���V-M����������D8`y��<�D�Z�5����`ҵ[���X8>�Q�+�Y�m�L�Cp5~"�i!����a�
���	�MO�����B�"��2�T7����\A�I�o�}8�àq�`_�K��w�.N��<�_��r+���>�m�0!��	�?���c]dkjd�9�f};OA���HGX��[[�klHR���B�I��N�-%=]�$X�v"ɑ4n�<���v�{Ы����1�����m��(�_?�'t_'s��n7�Z$qR-g�}�����
�3�U�	�ۉ�Bk��c�4Ƕa��?��d'L�_�� L'@\���P�>���u�y�f�O��1;arQ�	$|I�KՎ��^nKɳ�4X�,D�|��"93��"���$�7Y��y�������@�N�K�d�ct���}u-�D��g�w35_��e� �2ty���dM��E�Uಷ�'�;6>���X/�I��>�ѱ�*&��7_�~7$c[F�O-n"Y�'������N������-��C�*6g�uv�����'z
	��r�/@B����p�\j>l{� X��P���z8�&7/o_qq1��w�7~Gg� �5��O�|��Ijs$����md��41��=�Y���E"��ll�]��wӵ��x�aΗ�����b���w�{q��lO��5ޣL��3ZVZ*���L��6C2�\0��`�}�^,��J�t��B)��x�K��x������$zU׏׌<`ۋ��s�.���]�J��ˁ���#�9�!@'��q6���$�����/%e ��EM���ˤ�(r�1��zI"���� zZ�	�����߾=JM�>����WW�e��Y���9m[9L�(�������[��K���G---����f9�1{RYQ��&c�.E}9�]�Q���{K�r0?��%2�%�:^3�YO����?��dH�UND�k�@ �lz����S�9��Fp4�����h�]�|/�5�_DJT��'A�����^AW�H������ b^��z�����z��efeU��Z�D"��e�wI�o���Һ����%!��k�K��n�^������rs;k����W�+���Ȉʷ��o���MI���Z�]��󘻕���w�C������FF�@s�F�j��[�,�HZO+�qm�n���@_�w�{����f���w�_��6r^�@�I>pC*�ӱ���q;۞=�)�@e�A1�E#I���+k^.uK���'jM?f9� 8�� S�@�T��.��w�=��U]dnI�p���{��%���kS_���S'(,�Q	f��.�����f�kn|���Q�+#��
 ����g�T/�����Y�y:a�x�[�%���*����f�4UQ@!/�2��p����W'Xk����u��ӧ��e���[��S��7��c}:[w��1��rv6�b𾿫�a�g O^k8��<���f�\^c\�s0���Uv��w�
ܲp��V^w�� ��;��?ݨ���MC� �M:�M� C��},\K��RZ�B�&� xVZPp���X�{��E͎�Ύ���S~�=�y�tWj@�XV ���<G ���ؓ1�;Zv���5���Ά�V��l��&Z�	Jh�^��kd����o������������{珰���6�)���i�,w�&o�@�X$Pڡ�� �4���Fe�)<�8��O�!*7141	u/6U\�� +܉i.��0��O� ƺ�:w���f?^7�^,sp�f��t��lhf������8U /���@����l�T�	�5��it$�ޘ��%�O)>������Y{�h���t�����	�m�ja)P<͇]����(wY�o-yꔧ�Z���x�[�'���<��G(�mm��	��X�����Rp�[`)}�ROG�H��F�E�8�3�	]��}��m�L�Z��k}�ES]�w�hA�r�����C��ќ����.�&��-uC����|7˴{a֨��fvXq����Ps���<{�#S�Z@�S�d2����U�%V��ә������q��������^}Avֻ�s��j��A� ���f��U�(V_�N��j���3E:�SO(7�|0��5w���P\ؿ.,<�<g���� ��Fe)�X+H$���4����F_YLb2���D1�_ל��.
u�ԩH���gv/V�O*����w���AS'��EA����K�W�"i�Ts��_Zzz �XPP�'f�V�u���7��:EvQ��~��}]i�Z���{��oG�+��C�3�p��HF?v����;<=�Ez�����&[���j�����$]�A~~<N���ie."��Je���]m�=ɧ<���B��p[��k(���Z�g�_ou��Cj��Z�7�]��:�/EEhV�Y-6��L �W�u_�X��M���y��J��z�k��/-d�!B��������ۤ�3�6hBU��]��4�,��� ��%���^�B	���������6�F���ă{��lp�őhF��Øq��~�,�G	�k9-WvĢ��p�@SμL]��.�bU�T�99b���}8�u�HrDq����\��j*bcku�M#�� V��Rh ��qprR�z�"��ž�AQ��ĵj8�}}�EW�#���}l�<&�8�Q���xr�wR��`��Mӫ�
�A�M��(ƭ���M���o�������)+۞$�ƶ��J�%%E�]}SR�;j���oԦQx�])== &8�����)�J���u�rY�o	���Wy{��_�r ��Y��=�6�WC��U��<�f�i"% �k��3r�"�zC�����gC!�,�J��b�~�����������n�	�6tBHB}��z�����d;����8GRdg�w�c@��
��l�����0YeNl{JJJtqեӭ��d����(�ȧ�����tl�3�l��vd�gS��J��I3����?ͱ���6m�c
^S��IV=T���ODy��t_s�V
	�]���+�}!h͟;Iv�f�B]Gը} i���4">�)tf����<4��:��J�'e��-�([.��z��.r�)��M�o �0d����wHGܚ�/f��?�T������K���k�=�����o ���>D������C�5a�]���+y��_�������9�f��*�;ǃqX�U�^MO�p��L_�6�p��͆7S��> H���j�8}�N� �V�5���ւZ'��QH�������9����Lv{�M5���;�]:m��{X�yx6�
�U���ꦭD�X��l �@�T�D�)�]��<*la�PWo���ux�j��rF��!�Ne^p����O�̸�t����_�YC	R4���&���JJx�Y�.E�ɣ��S���p�j�T4�J���қ����g��.�Q�'���E�'�Ν;WF�삭Q�f�j���1�6���ک�<�éQ� �e$��ݟ	Z�Ys3��@%�-bz:T�)^�/��~q��SfK%�/��^6�ʯ�$�DY��� �O�5쳳�SF^Wm�+$Q��\n�$ �k��#؞������,��I�#����@+p�J�Ȭ�>����"̎'�~�����o�ċ����GX;]�z�@�~���&_֟˝F�49��Tzϒ�V�����Y��s�3�g��`,�H���k��yl�=���9>�745M����j��Ry��w�TB�M��	~�[� ;��`�h<Zg��~�v/wu�4����6Sz���J�$�ZҕђH]�t	�訥#P�>]�?K�����V�Q�;-���RampX�Ř_ާ<Q�hߤr���R��t�lΣ��D�Pܪ�=劲�|�������e�]��cl��֯�R`�,}�6]���.��Wf��\+x�+��W���s�Sk��q,���Xwi�Fc���}Y���l(��+��O$.i2P9ި��҉0r���#�h���ȁ��co�M�͡O�0)�J�[��� �������𝮟���S0x��1�a�tB9Ɛ�`�G B�KT��Z�� ����d�|I�u��]jDؿ���*@���v;�i�U�2<T�}�rjk�e��i��������Q�+Aw�&�e��=|2;�����R\Z]�:�$��@�%�1�z۸YV�(P����Ŋ��],�|M�G"*��q�j��r�J��,y�k��䐐?�#������������&Y�]^U���3�8^DO,y�w��\����>V�<߱���(�@�ƠQI�k�,�س,//����,?%��1��˫h�g����Է�S�Q:b���n�s�{�wͼ\h|�"���I��)�i��+D츷��� w�Ә�i���kÈu��u`�����$���v���-T��T,��UE�K�X�Q���g�P�A�fؙw��a2@_��5��8�'�fyՅ� �"����ay]>�H��'���$��[��
&�Z��}��*!Hu!�s�x�h(��ݾ��. h�P�s�*?��_�u��Nm�ݝ�~�C�V����������W5S���7�x�L��h��TE�|�A�����A�#���'��ݓ4[6�Uno�vB09;���L����;��q����d�I�H^�77��7o�G�z����O~Lf]g��&+�k%}pM|$��KM�'c�Ck��Z)G��B��Nii�E��ih~X��|�~v�l�r�M�����J�p�sM����bta��I*���f�����\W��,�c+$M���g���Lk���6;Zq��ɓ�c��m'&&X��o��[�VL.��dc�)-���%���w<���n:���R��l��H�cW��)�M=5��KA8�{��Lj��r���s���$�}a�֜_�  �S�O��w��>�ɂ��B��������5R�Ua0B��[�2���Qq�9�#�o߾eZBlL��o����/ �����������X����gO�?�7���_6����j����H	�xr�M¹�-g����3�ƿ1(ZӨ��i�#�X��IYQi��(�@+h�X~����pG��E��֚�(TU[�ԂH�}���S�F^��<?k�PEU"=[+~�C#,�\����RqQ�M�\�O�0�
){Z�5_������֞���V�i��mvv��	��bd^��I�ø{n�x�|��333:P�����A�p����x(ӎ�����AqmN;UO��	j?p���|`�g����� 5aW����'?p��%o�
MB��ϣ}�`FisؾȚ�7����nM�brA�
�	���/t�2¼}��Y�0a}$cIS�o��t��R�A�(�6���:��� �<J;�d�X�bB�xZ�ܜ�_�OhP���=�oI$-�p1���-��'� �"�(�U�	]����^��9hbs����ؐԶb��:%�ؖ܅?���A�TS"�n�i�'
�P76+=�-GRr��fjs�U$�~0�&��X ��KӻZ�>h �q@�=������J�λ:�A	����
b�<� ���ݹ�_[|�E�jf�)I>��� ���U�h	$?qq������\$�[�W�3!�d�&<f����Ļ!������~qm ��6|���TLX)���<��Ьw�?�-�x� �1 ��!_���C�p�r�~�M})�y8�7� ���;;;i7����h���(TPAHK?��꿇+�U:�|R�(��
>8?]'˞Kwu�12�~��Bo�m�C�O`i�;��@��:نJ�V���#1�!����>��2wfD��t���^��s���0"�Wh���[�m��W���-��!�`��gc����ŝB! ��84s�*��IQ��@��8Ȝ�995iz�� ج��\ޒ1��o``u���o�><���[�hȽ�����M�v�@Un+|��Ǟe��� l5�ѱ1���k���aY��T78VFy�����/n��R"�k߹s�#Z4�4�R���c[^t�BF�wS|�#I�n��Ѻ�)
u���T'S�6����w�0� �����/��h�>nAd������?mP�}���M���㝅�@F��&���{{���e	���Yb�����A96�	��='kYq߶נ�2��7��(|]�_��J5	�Om�����r�;G�����fF�6�]��+֘��}�H`����у������O��(t�?���̗���vh�
��2��/��
Ƚ���p�߫�NG਴CU ���{"��`������z��7\&;{(�t�u��V���D��+�n��SRI��R����n��}��V�翐�����2gA���r_:p��(� h���A�@�5T��.�4Y�St_��k�ׯ�����`	���F�s=S�a@_���ͧl�����9�k�f
�{2��Z)pڄ�"�<�ޅ>����% A�
��i�t��rmSu���QI8c0TT���w�}g�w�燼*�
��]MG�A�(�q�F��IԂv�<'��y�%l5���l���b�V_�P'�K&��!r�^��%�}�i�}�=%2���Ջ]{_dgqx�>/���TF��=���+��z��h�s�n���w
��B���u�:dt�P��x:����ms9�k!�t��Y��n���c�p��ۭ���T�is�-���R���w�@mԶ=�_V\�x#�[�-����������`�ݸg����@�b˵- a���}1v�bon[�]��_���&, �b�a�7�I �Љ��	� ����
����䓟�1j A7Q�Y���F���Q�(рN����goG//L�a��� �,�g���:8�uX��7����{9x[�?<�z�>�/~�s<�?��m���Y]�5�/L��<�ǲ��o��oT���u��������޶G�8K�6�.�f�l�W���t��Z�~���~�F�����ȝj!�FQVgdo�S�(��(���y����e�D}z�CдI��Kg�˶�I��k���/�������ہ���@���o��ÓǠ�`y���
����}y-nVm[qLbM�����A&)�9����I�������.4�՝��WĦD�BzDm���5�֗�.�k�����z�e�� Ɲ튌)(2����5�#=@���S���hZ0C�O2VO#�n���K;�T����\�r�޼��w�rq���Ѭ��e�D[�+�ڶ����qO"M�-<�}���L���]��ҷٗ�SH��^��ČG�2�	�+[��H���7���2��;���S�mn���4�͛�O �a����.<���8�~�g����gB���	�׹�N������oR����,L����O��Z�4{��/�%on���3��E��Yږ������:�z� xݼc�Ti���%���JܰR g̚@"=�o0IB�b6l�켖A� �8�z�#L<ՈY�:ѹc�aa��@\˨�V�{m���n#V��x��>���<K��au�h����d�gu�;u����8߆y^�"��@�`���T�1;wI�/Ok���B�Dܐ�����_F�z�!M.��u��K���r�%��OV�Ն�*���	^��~�sbp��&Ӊ�i�B^Se�}�q ������[���81�ǘ�DM�"�D�w��Sp���G��D��D�����)��4�T�����::2z��� �1/yN��1i���3�1��!�!�?"񗈤��}8o�5����5(1H�(��f�����K�:���r�W%��TWDۋG�(��^g��º95�dro�N�Ж
�
��D����!_语z�X~�F�p"�^�h4;z"�&52I��������F#%[ \��Ng&uY�u	3��UR������j�Cʴ����kJ���5�Zn�W���O��T\w�B~s[��r��h�&l���U0�ъ���������u=����(�W����FVrp���o��M�f�-��{_�:/�K*	��	׺�l��&C灧�������}�����*���j*�uը��ΟF��1�_0li������O��2B���U�e�St|��_�m�+��;/�N���L�X0���U{�ét�V�Kx��,|��/Q���W������NiV���)��;�TV$&X�q_gʗ��Hʝ�~���{68/'�^��������RC~���p�LnE�����bt�%���qF*Ӎ��Z�EK'�7�\<-ֻ@��ef(vu��ZYmyB�'_���Ǵ�3C�n�S�O��J�H�g�B4����,�����n��ު҉���[� �=2�&�mU��}�����_%�)��	��U�;����3�qY��d�OUg*�?:o�\S��w*9�Zx~ �q3������%��r�if�W�x��*o���R��	!���)7�/�R����Z�vJ�az��a��V���H��A�\�~��Y��vإ!<ĳ_wΡN%f�W2�>�2����P8���`��o0�'a��_3f�P�h:W�6�	�(�k�2v@5�?�4��pd�!���X�����VB�̡���&U��Eդ�(2S�?�McPi�U�2����5;|���&�-�P�њ����+�����4E\������//	o�+�Ӕ7-xj ��_B�*��f�/�;�yd"y�S���Ā������1�q�ܚ<<��Z]ɧJNm��ޯG��9�1 �I��i���U����y+���Y�j�;����307MU����#�(юYK�����vO�h�x�S!񥘘��~��WGK����>
��$���m%�JB�҅x9��f�g�%�iz���8��-���b���fi�����u˯'Ȇ�/7=�ߤG��i��؊I���6��ϴ]jiӸ�s�_�ߌ�Q+��<3���8sO��ȧ�ZR�7\���q�c��*q���sZ�����G�_O!����5~�z�Q;)w8y��Hd��O�o� ��9�S��&�v�`^�� ���q���	�#�m淪��[�>�4ɼ�(�$PwA���� &�<H���rƌK���$� ��.zJ�C�G�m�߿/�3S&�o����^Xs�>�t�k#�}V/�\n5����X�蛺4��)���+�:�6���������¢':7����蝈W&������H��ԒK�E��R������ϻ�8��\W_�;Ж?�������;��[�B�ԩ�)�Z���R#_�g(��dgg����S·"�O�i��vE���o�����!1�1 ����k�_#����{)w��-!W^J� \�#��#�EEýK��i�=��/]���xxh������i����[`糼�^�o�0�LMIe��Q���G"��ej�I�:��j�$�]ۓ���QQ9~\�i���8,6q����GDD�p@�Ѯ�Vz���сJ�c't�U�ȫ�Ȋ���ݽ�|�U�ik�x�u��]XEj����&�ʡ!���P5���p��+R���ے��(�e�Z4�@c��.���D~e�q�#պ��N��>!���n-�șH��<:�C�rr��� Ä���_�E��'�L22��<�>>>Z�� �A�a�X~�b�S~J��z�~�E��L��-��&V{�Aȧ&����Ԅ�W�����.���_��4d���zx�ė�i�ɬE$�D�듹yմ��x�z"惤
�4 =dm'Iihjj�^��L"���T���nH���{%a�T`9�O�R��7Z^u=�U�+db��C
����A��6NJ��=����)4,,J;�}�[yn�۾���p��U%^�Hq��CPV������OR$��mR����o��`���JC��-�H�u�B+F��Ç6��ꁷ=x� �,u@�L������ᝃ%�vmc����c���O%8t���������^?�����کS��[>
y�F��25���hW�ҁ�&
�^��lfC@Ǐ���W��;�|H��ڝ1Q|V?ʳ�q����9^899���Q�U��}�����2��3���v�^~(����&���j���v��ỒWJ�l���)�cv��L�>���H(.X}$w8�������`"$�B��#w@(��k>�cZw-��"k�����bm�%h]�E��)����ۿ�ل+�У��ī��-4����5I�Y��tx�+^'ܔԜ�4S%4�5
����l���U-i| �L�����ӻ��[�|0�	���c����\v���ml������3N�_��Tg�H�UY=����4E*��������i{.^FZzom�dHYY켃k�<��v*�~F8m�W�9�4���1��o%9AϿ/��z�Ds8g��,<���z���4�A*�v�!P��}A�!2�Ǥ�`)s>�7�����W/N�ʥ�:��`�5Oԇ��ntGC������^����T�������C�����R/�@�o&��k�B��7
��D�7��[�tᲄ�)䬧�|�����7^5���Q��L�ʕ+�==��TL>0Og��+5�6B����̺���3��.M�ូk��ϯe	?��9O�o�f�7��j�MҎI��sc!��ă�+���/�<9�~�5�+y�ٝO��3�[;ᮊ٘�j6��~�o����W-ws-��E� v?�[e�|���B~:�~8,��*mM2���j��Cg�(\��H?i�C�v\�+
�#���xEnX /@���-����W]Ԧ������ˊg4����?đ]��=�{+7:��z/�Fr��3�>��@m�����ſ��E�eu�9^4��l���V'��s,[i@ἆ��@������"�B��?<||��fR	2��+[���Ow �pRj��w0_�m+�vu�-+�i�2W������ye�z��g��Ď�I��KO~���a��WJ�yp��Ԩo�Y1��`��%2��Ǿߴs�=�>(�"�	���o��ci ށ;!m�.�J��e1�oAߪh��0������a)�.�}���I|`�(X��8��EO���&�0zéVׄs����gϞ�
>Ua>�g���;���VU�����M��BӃ�!D���7wj-�����9�K[Թ;�U^�	+� _�q�X�AX���\Y�mydW���o<ԏ�>�}�z�jk����-�!�6
5$�ғ�T�1�8����"��pE��Ґ�`��eW�W����ŋ]*�5Ր��iqB�T�2��=���f��iiJ���z����&#���/���[��t�8��M��h���#4����Bv1�py�85�����j�Qe�ѹ���t��FE6q��^%S#����56==���S!��M]ş�Պ)ȝ0�k�B�Wͥi��2�u�`J�篢���w�J0S0�Ƙ8]�gnT"a2vy���>�q�{u��f� 0�|Z�ݠ�k���0�R]أå����������N�i�c] �02�	o�./���q�i���ʒa��4悙J
�Sh{�b�l�Tr�5�����dIř�W]�����bk�@i��4_͵��+|�{_�bֿ�ߑ� ��jqj��[Q�K+s��AE�M,�E���Gj#\<����0���dM��ORV�bJndE[U�����<z�h�A�/@&�~B�[Va�X�>�n�mE	�����:w� ����d����:.��C�K�:t���K0�����3k*I������Q$��󱀹<���V���R٥sm_)Xl<���QU��^Ԏ�� R^�,g�[���9���,�J�YU#�b���I�dA�;k؜UDh���F����<3�<��6�;�G���n��$`F11�**��d9�%랼#��X4���f�;��86��4�IE�A�to�����k��"�4�	�E#X&S �T��鈂�j�����j��h���¹6����� ��	�B�.O�-�DpܕY淼�/�����߅�' o���h!�A�|������O����m�h����v���1�l�I�72�m�ւr��� ���A�4q�vg���/e��?@�k,�ȵӻ�����A���3Q�w�Ų��	A����3�{yL�5zE�������rT�����/Y�}>��fZ	����\bW��6ߦ��ʷݎ&˙({Ǒ�H)�>�'@|6����a��E���Ϲ�X|�AW�m`n[���;��Ż̶��|��S�Ar;�Sr�
coǼo����щ��]X����og)ͦ-�8a��O
҈ޫ��g�����|eN�K��%��ǽsg��P3uB�����V'H3uqg��&.� S������P�b��%�M(�P�#R:��m�"��j�I�<WU���d�WWpŃ�-���ϗ��r�\ANU�Gw'M֦����}�c�O w1+A�m{��ܨ�dNz��D��D;j�|�?�����$/:��4�d���������QN�ϴ���Dp�FJL̆mJ��׃~�����5�ة�RN���
����A��j�F���A�e�epϘ5�H{!����]�����"�&z!��#�1�/��ѲL����k}�F����KJ��'�K�c.,�\ ��'X��>@|�Jy-P����q��BG?���(\�j+o)��,�㥩G�LL���qI���1���t�9B�%�Js55c���V�<K�R��H�"o��E��B��zsZG �7r=P��~Y5d�eU�Ĩ���G!�i��P�J9;�7-^.	K�Vݲ���g���[=A+v����|ױ�A�7�o
K<iw����:'''@����4+%����U�h�
�n�T�?O:)��U�-�}XT�Ջ���4i�_�}�k�$M���2J���i~�KX��Ț��$Kޯ�$�H��t��+[�"��O���r�xaԾ�����M� �h�H�'�,KF}�Ň�|��kj��+F�í\oV��+���g��8��(W[9.w�^�5�Dݝ|�ar�y�}M���Fg�E��C��ے�S��.�����ch٬dNNN~@h"{�ы�؃!���e%��_++}��$`���i�J&��t���.�4���_X����vZNR�>y1�iL�!T$^w�'��S���\	u��ŉ�!ϘZtG�4b����Ȉ9�;Ӥ���Ғ�J�w� ed�y���a��9=zd2���ZZ�6KԠ�H�{#�I���T?98.)D�����J�s��sj�����{��.Ȋ�W*�.w,����/���A����B���͜Mjƃx�*M�F�4�.���냺vtl�@�'IY�B��
fw�u�neC�X�:V��wv1���쵻������G9��W=A�M��q��-F�N4��������Y�ң��VSID�)@v��}�+x��F�}��=Jfe�1�.�3��,�^�tu��#��w~R`�W�WAAA����Š�ڬ�� �R�vQ�]	T����6K�Ɉ�-T�$/��<�]�Z�ዬn��IY�?2�����!B��e����<��RDc}��0�)���볁	����>͔H�z����݈׋u������n�(T:q��C4�uh�:�CʩM�u���\��.����g��"��U�!(�����Vۣ��0u�L��Or��Ԡ����~(��E�]��>?�i_��r�k�w_����(F�.6�t����'��(k�X|�o��꣹��A/d1��b��qMh�԰�ǡ�
�\��#N_�?չCR� �E~s�2U��"wl���E�+�_��Nl{�����s(��<:���2W��l����<�rW)�8���D+V��*����Y�� ����v;!1:�0a}�؀�X�|��U{��n��k�j��XYN�p�oO�.��EZ����]�B�ռ���uv��&�3d�5��+�����\��{��*�WEn?V���d��k�8x/U��@r���>Wo��@�ӊ=!"�ǫ���o�"/��(ned���7.766�&5]6�d~X����Y�ߗ/���m���c"9o��d��"�1(�A4�= 2� "E~m����ņ2��AYM�OX!�u����Hƹ��e�Ӈ��V�q��7�1�m��W�hD�+��B�=tas	����Z+��l\D>��-#�=o���*�0jݏ�W���_�]nr#��RQbce�c���Y ���\�:�eu�ۄ���?$ٹ��?��w�Q�0K^�L,&�e���%�n&�7�&����f|X|/��I�����1�sf�x�?�v�Ӈ�m	�e����~���@�/���$���Cm�6�G3��Q5Z�n��� c���������F��V)�Ŏ��Ģ�����9��bE"���k�j&�w��cO�K�1��W�'�N�}HSUw��I��|�%z"ᬱ���_:���u$U�Å;�(V�~�Nh;l�X��Ԑ��P�F�YxΉ���S��.~��*��	Ct�8�2��s�X.j��:�^��2E:aO���R����a�T��Lw'|�"�l�i���gɵ�x��'ѣ�6��FW͜qd�F�i��������x"2�5+Wh�u���Be����I�t����9�VkjMt'��V�`�(�@ݻ��#D�:�C	�4�
�:���=4�N$T�>;�;	O�����)0�>r�����+B�!�ETz�gS5����)/$P	��&��d�;.?�;�B�� �^�_˲anL��)R{�[,�+5��g�..
wSn}w5F����9�:���u�q�%��SV��Yw� �,b1P0���r%7�&�I��5F�uZ\W�����6u���3���4+�76��,�p��O�C�H�x�V��[�>0?sz�Ze8� S�l�jh�v�@"U�Xw�����S�Q����g{a=/�}���É��R���=Δ�/\�g>�`�s����Y �_���.���氂>L�ý�r|~O������d����Uo���]�+E`��E��@oյ��gJ�@��F��g��!�BWz��L��m:�6�~�I���
q�H�.]���y�ń��v���N�����y�� ���/L�0}`� qD%z��,�r|RG�\pĖ7���yN��L��˴J�T�ӝ���)�o^S_F�j6�����$�OƎ�B�~$��E����a2";��T˓�,�-��I�Gx�b���i��1U[�d@~*��Ŷ�wM��gU"�o
����T%�O���F$���	������y����'���e�|
^�߱@������k0/x#<�g�}�O;!����3���e�0r�I-"���/��Ί�3�>M�֌��>��r�,�;E���O�^� J��!�m�mï��Ὧi���䊹���W����RԽ�r���/�%��^�d���v���K4�w�n���Ga�wX��dH,Tt=u��O-_Uץ�����5v�l�.ߐ��X�u#{UF�Y��1t��'럯���:�T��ax6Y����!��Q~�`�	�1�٣>�m�Ŝ���j{;>�
Ψ(�;g�Q���t��D�^"n�2�V�}��1 ��Y��VU��a�yNJ��(ލ7��V���5`o�����_Ƚ��Ӻ Ü�rk�0f���Mp�ծ��U��2 ���jK�+?|HIo�21�G`� �5��}�Ŀ(J~1��I�m����V��j7g��rY�|2�M�s4E/����#�/���8&�4�h�|�xV	;0<�e��4t^H#����Ǥ�)zƫ�ٹ'Rˎ��o��!D�T�����_y��S��&^ܶ#д�%�꛻��7;^�`�V�z0Vy9^�6�uou�rj�]"�(�8�V�V؇�1��������}!�s2l$�,���ů�x���}%q%�zl���*�qg�>vr&�i��[��5���_|ഉ1��U��&��ZϠ��� :2U_?��� -���	N�{���ݯ>��?���'��~Ǫ��'���A����E+S�ޑ��#�+�)0{yJ�n��%z����8�����x@�p+��ƿ˹\����8p쎎6��^4�F'�w�cO9Į^�cr�%J����^�~��vz.{:��f��9�St�J
���#Le�G��H�6z=n1��o�`W��+o�g��"�<���F�[��;:?U�� �˒�|��SRxv�y�Ԭl\R�AJj���nN���(rPG`ަ4��p�ʤ0h0��px�6��§�`r�u�����mv�N=����O~�)r���e,����.a�����O�/���W����m�@��3K�W]-١»�$��ړ��$r�nm��B<��k���'f�إ&���jx`&�_�R	݅ ��٬`�p�C?��=T�=*��$��.Fk�"��#
tJso�?9�j�y~\��YX>mR�i(�ab�A��� �~�����C��9,\�t�)���>+bƺ�F0R��$���+q �����Ҡ�!
��6U��i���vI��Cv,L�RlU�EK���X�e�o_A�~�>6�ŏH �Ib(qTrI�ɶ�FX��IR�\�u�|�x�ͥɁj�1�-�a����h:��������,k��AP!TwUP�"]QP@Z��J��KG�zD� A:�C�	=@(�|��Ͻ�����������9s�甙9S҄�{�|e�A %v��=3'<�9U�ԒN|ќ�nM��XbہK�ڃ��,�ӑ
�w<7�6�׮�K�~��-��g�v�Ս]0fgVQ.��{U��yt.� � �w�v�h7u��R�9�?!�:M�=Q]k���ء��;��� �(�� LYP%k�|g=>J�ܳ�S�0�a��8>���p.��=�õ�#ůY����Z%6�F�Y#΂�Ne����<����u��S��L�nt����5�D}݂Șm��Ր��x�{a�r�ܿ�V�x�ᖅ/�v�J�]����h���bz{�Ҿ��E����
o/i��������H���k�;�}Иn�Z�oN�����8Y6��9u��=�W��c�ly�ӎ<ǀr���3~0:^{��Pm���g��=����Q^XF�.W�����~��ǈk�+�aG�8֒}hkMT��s�w_�MI��m�VaQ)z+x7�Oo��Pl��q�O��W��6�ї�)|V����a=�l�Pva
��L�-q�#��)�{R0\�@y�Yb�0x�u�E�/�i�#i�|�k�b��tJI%�RC�?w�^Xn8��|*������'�-�?�e�9<�fR$4�V����<������y �Q�%@�q�Y�'�k�d�W64[<����ɡM�eȺ|�r�E��V��W>%e���y�:yczcF4�����.j}������n�31}5�,�X�d#���
�!P���+o����ہt_:音=�]68E��ˌ()�������<Fw�^�8.o�5��:7ݙ������K���LuV�_@x�����{��M��aj��⮶��m�2_lG]�)
�(��	�ˆ�alR��#r8�:S��%)?:s Ko|�60�m�۟-��w$��b�#:K�M�MIzs���BӡBߵ���=p?�N��`����� ���8H��j������~$IX�n�\<[���}U)CX�'��e}4T�Ua$��@��I��mo�M?�W�Ś����Wjn6'������IԄ��FX���f2�vY��>z=-C�ֿ�hH�I���;���P�:� ���n��Y���ys���7cx���t�E?/H<	�P=_M$)bR�����HC_J#wZX���SPJ㨚�a�v�!\t�"C�ѩ`�t���3.S��+��!�}1ݻ�m������lA�g����O��*Y��Vj.��M�I���P��R�;�hv��a�f���qC@9[�3����?_�����)�O�B���2�-�b{��V:��P�g��a������� 	��"��7�F�ﵣ%���_��%-�</�s��X�әU����K �����8���A�J�Ջ%6j��T�R;�]���}�겂�<*��[��I��sk�U 2z��v�7G�q%H;��(	V��K:}zEtRoo��8y�;�Bi*�(I��g���w��/�]��~Bۖ�f�ҞD���G0=�&�[�.)u�"�.c� ^�����$�i��@j�M���)_KP0�gl\g���iEԶ���<��9q�w�R����'߶;��k�bt>T�y�|"Q��8�B��E]���9f�ze���4��V�)�#V�Ћa}b����(��.?|b����A�ɬ��ԑ�%r�
�(�lUGR/�E9��.ٚ��y��`LdfNE�`��>��RV�>�U�M�p��M�X<�j �Y�)���6���o�&�0#J��F�MS�eE��K����4.�g|"099y���%[I�RY1";u�'�}ݬOW��nʤ#��})6���,��V���>S�K.�k��Зn��􆧚q^��.sX�qFb��p��~L9R��3H����k|�m�<�N҇j�jSw�l��Y�:��-!�gn�����m��E��_hL�Q?Nv,�k�M�!���]��=JT�w�?~����~�Ѝ�dy��*_�����2��v��-t���Cw���V>��R�^�a(VD�4�Z��]H`@23�p=�v\I��
�._��JܸW���γ)�����i���b\cLL�P�m�����=9��X�
��E6v[me<)M@J�^��Q\�ѣ� ��~~���ZL��5�؂N�ϘN����-+<�b����l̢B�{�K�;)ʊ����|�ϗ�{{{ێr�!�h�u~t��1�.�9̖p�y�ISt�)y�Ҥ�ECc#2&��C�10��{�j�ڠ��_AW���rx�0~-PIF�L-ʊ���~ඨizL�J��O��߄y�e�~�|�ZDv��*�%�:n�Z=v�.�-Mb��!6=�ĥ��g�2��vٕ��v�����Z�U��T�E��^��gWl�{�J-�s�����"�Ss�,����ﰌ��mD��aiR{�����N�T���-$xת K��z�R�Я�_O�×	����XI��HF�y�=)Ob�
Q��UJy��<�*���G�N�K����Y����j7!�R����V��0�;v�x�R���T [�`���d.	���P�fj��]�c߭��?��,V���������,g�lҚ�(���˲
1�mé@)�'�:/tf��z��ݼ�������̃�qq+Þ���������(���j����{
R1s|m+��a� :�<f�Nuܮ����!�Df�"8���W���~'��a� 6�ˇ����~�+��B5�Y�u�nP��ľ���N���(����OjM�I�9G�@ny���&�`
)�j6N� bj���t�]|u�E�L~+M?�l�%'w�b�'@SRT̗� (�h����*���������;2 `����zj� * d�v�i11��:�u������'��6%%'�*�d��\X�Y)�S��V���~�\3���"���@0� ��mT�d)����;G��TTT�f{r�w(�>�<6���c�$�e-4�!��e�j�u����u�]�����Ri�-�����1---�E˿1��z!4�mj�>'��6� w�yH:|] B ��(����4��~'��;� %�u�
�	;�"�1򷳧�[�s
��iy{���B�ҕo�k-PY!O#��l �-H�2�ӵS�S@4q��an�KP%����2N� �̚��Ó!��7��Eށg]��3՜�Iq~υ�~ ��	X,�y�Ɨ���@����]v#�������_��� �}��J�j+z�}ez�ʂN�a/�$$�iX}�O�w����d�Ӣ�dM����r �Gc8��ٯ!��.�����_��	�Ċk<�Hŀ�7���5�%P��,�ɒ�~��nw�y,GQ�^f����ߎw1-mhԎ]�z��`@R*�Ĳ]�E�	8z�x�I�w��X�S���o�j�:�gg�n��o���
�6,�ˉ#�ހNr�~�E ����t�t�����U������\��"xSy���� ��q8������v7�����I�A
P�/��-���N�ϱƗ�rp�q ���#K� U�������m��{<d�o�h� ݪܴ�yW��~a�:d}> ��v��@p�5yZwY]��1�m44{�l��a���i�D
��ޞ����iu�҂���֌1�;��-d�
f��t��n�o�W��ٞ���)�)j��$��{ZZV����Q����Q�ee��s�v����ͽMH���אZ)0��s;�L�4��&�ᄄ7D��9�IK�����(Ah�7��HڏݎE8����}�^33775������	��V�����t�?���n��.J��`�1����� ��m(�ܞ������FUM(�{�!�x'KP�����k�#��~�T<��Ú6��F�d���~��	ĊW1*���Ħ���X(�.�HC)�E��c����\��8M��A5�w��FgO=��dTP��6m�2���/(n4]�����LI鴨	�U��&�]BA9��ʏ:^�A�O������/�Q�8b+�vnJ��K�2���������2�Sɡ��8�BP ��2�#0� /��h��j��>���SIzJe��՘fh����/���اW��z�"���N�+��?C�+�m��b�9 ED7�G�H\��(�6F��7�ܦ�����v�C�Pi��|�d s-��a�r�E�C�\��ֻO]�����/d���n<謥���*����K�$e����Z��%\���6AqǾq�G!t�!��yw�	�|�Wfd�S�<��9q+4�N���f�MFW�G�:�?�T�}k��u{�4�8'��� ����J�&
&�=ؕ`��9yy���S�n@A����G�Sz���8G�Yo�ԫf�h��@��h�kV=��_��UH�'��r�H��I�s<k�lKb�:��	��(V��CG��b� ������k5X��J9�?����JA� �*~@U��0.{�0{4�}�h2)Z+��t�ڻ�C��淎�yQ�2���p5p#��h�����ڞ�.�Az��
�#$��j�`ٮ�DC�+�޲�v9%�<�H��S���Cϡ��8-��Ժ�U2�nh���e��
+�P�9 �@�߃Hw ��{�@�����d�׾s gM��R @&� �A�nfvncc���!�)�]�����B����xf�Ũ)T#nGq��)�:zX�[Q��η��s���x^FFF� <�B�y�j�uc��^�����`�ߏ��u�W�X�S#E}��4G�>4feʧ]'=�����fv��q���2 �����r:�
�������@��2#�p9�W��C��@�wx�⏸ot�B9�ͣ��}�[�P����d�V?($1�Z��ʖR����p�ii��ܦ�2�g:��`�F,�ɪr�O�Rq��7�Z����9;(*� �5�-]ޑP��Pf��>"Pu�-4""BY [������8�TB���Y4��|h�֮���ܮ	��Šѭ�:z�ijiힽ���bfީ�mM���+�r��kK��T��A�y����J��zKo�R}�^^.��]�NS���O������F��*���f(�� ,��9f׿%<� �VXq��2.�M��^%F�-F�k��q� ܍K�t|���S���q=#ʉ5e����h�*����p�w�d[�-B�$	<���w�j��:�m_]cȟ�4uɱM1vhҘ:Ek������L5N��8�CqL뾄�ⓢ--�X%�`׻/ْ.���,�����S���`�ssj5���T3h����@_d��r1��'���/Z���Ũ�S��ܵ>��r������D3��]ŭd�����rp�n�S����"bg�h�U8ݮ�͒` �*/kl7 �_���7ٿ8N�����H|��:��Y��<p�E�h��Q�}���<�)O)����f���/��W�rpqz��芦|�f ��M�_�e#�s���0=p9�ec�4�<��H��}	C��nv�ck�@��;��8��- ����Ui: 3�|�hi5cLķuw�̓G�@xe��9 N3�H�.]���/���Y�?�H� ��p��Z�IEx�Z�0-?~��������a���i��1�?�D��WK�b�+7
[]{�f`N�����r2e��!�/��P�w�Ö'v8�5}[>tmt�V�i�ss(�x�N�|u���/�"5����#�u�N%��;���Ϝ����`iD;?�t�d������Rk{&U"����{���TP�k��[<����^������D����lJ����'Ų�Ϋ$�y
�U|�H�M���.V_�,B��.[H�s��X�l����g�6�����q�'��`aM���?U��ۊk߮<U7^ih�'�Ғ�0�p��_=R�kz���x�"��Qtn���ץ� r!̟M�[ګ�2�Cc����"z��������W�/ˌ"4o�ꗾ��]��&���k6겭�}�@��,�@��Sd�4��8�����m��zM�Ym2u����9����>��������Wer�Z�I�T��/�V�f��7i�C�-qdKf(m�j��0wf>���-�sಜQ)]w�.�Ħ����t{5�k_����Z��R��;�8�j{{Q�W}���a���ո����&{ٛ�`u>j��R��$����FX�����B�\9!O�?GW�V�g$�Ό%�oW�7�M����V&�_���P��A�窹�KWsf���K֤�p{�-�$
I��7����Pd��_�g^�J�\c���|ܒ��#�	'���+�B�0�}z\�*(D�m���nSg*�KǿMn�h��4t�����Z��yL>U����+�1�zx��uS�ZQ�!���Bq25�@!��v�>Fjj�� �5|L��mT���J�[O�' diҤxQN��\<�̙��E�G��q��������V�Ul���/y-�3���(Mk�Lq�M�G��yjx�s4�D�J���P^���@&�ңfF�މ~�s�����sJ�ǂ�mmtL��#�褠K�H���W�=����e�]�&$W_�����R&�ۑ���%�q�N(@z;&�`�3�[��n�3>��I���An�����VBԭ���S�#���j���}y�2���Ѭ}R�@;-_L��/���K�סg���{R&�?����DFW�p�����-r�E�5N7��'����\F�	���~cܒ妮�H:��k��s?�}�+1�<Y`��*�[��^�?0�X~i۲���)��>�]��������7�%h��r@��d����jbέΥ+G��[�o�_ q]���Cȁ�������!�QZ�pi�������Դe�Կ;u�+3�Wዑ}��ܥ�B�p����fmog��d��|���v���c!W�
��[��ǣ�"�Cy��ff�)������h����J�ϥ�#�[R)1)lpq8Gu)s-9v4 Y_��l�xj>p�Le�1���Ӽ(���EֆS�&��Xڵ�B(��kے<�e�cM�cw�X=<�5�S첤��Ի�bn�����O���l�)\���0ԨR�LگC���"�/) O�p_-���|�.aHnً]4�a�{�7x�D	�xb�܌���� �)��R��d�I궃R�B	��>PF��Z_^|3���������'*W�8e�h2�@����F�����te��/�{�}Ie�4eU�v��mll,3.��]fI֔�R�b\>ݭ��$x%ELJ��[-læ��+�HI�-���34�f����=S��Q5�QS��twN�sc���~tl�������7�N��4����N�u4���z������T�����^����;ȁM�`wc�k�m-�mx�&1�����Q����35����2���b���JA�� Cp[[*�T;|��4py;j_l�o}��b��B���e'�������)ug(y�l|o�[uOᩀ�[c,�rB�kn�/�O��i����%�G%j1�}������������L�%]�!9WB����5?_W͛���}ɺ���R2�;7����P�©�h��R��9�b����^ܤS��@�A��8�fi<,]����XNv�Y𝿐O)������P�	nA��LW��[�uF��ud��W����\p�"��� �G.'\�,&)3�ť�U��	O�隭�W3W|��!��q'�SiZj�0�d.��(Q@�J=X�+��lP���5�
\�u�#��ta�Tfwi(/��R����v�K8�b`�9�@�_��Y��z����E��������7�ٝ9Z=�m�bśT��#k�7��3V��XY}Y*�j,e�Rڏ�plC�����]����>���z���Pk�x��t::��b�ht�\_Q]	!���d��{Q^�����[O|^D��`����ތ��\<L�/��c�L�Zx���T5K��+#����Yg5�ð�F�&��=��.��%����וڛDb��]���9��6A!k[�KF�������aכc��[�q}��	=j��E"��aN˼+����y�D^��+J:��D"
��F6f�A�1�2��E�Ǻ%0`���FT�/��P&�]g�F-F
���fL+����}�����J���)��6B��ySݞ��,���*�0D�E�uԈ�r293���m)R���̠�3���>E}�H�N4ǘZY	w�����30C?����%�b��������i`���	;M~s�ŭ�g�Z�ϟ��4��Ͻ�_tp.ɿ���'���6vI�n��<�+��v�ߝ`��;�+�A�l�纇?�f�N	�K1+���;���q�^cZB�= ��k��Qʂ5*F�!km6>�t�\�Zy�6	���`��۾�����繐R��W&A��VT��2��w��c��b�2�m����ks#��wV��x�M��`�'Rja8e�@�W�����Ny�-xY����y8�,!�L��uj�8,'��uL��B>�^�Ⱥ�!�/�d��?����Ny�0,�5P���@��`P�������> }�=iǌ�uIS$RP�~Q�n�G��s$'�n<pxOE��R�$7�h�8��4Z5CV�Sjҍ����.���i��^�3�~�k�6k����Kͷ�y޸��@2WV�|��9�g���$
�s+��_%e��o͚�Te�
_����
�j_�Mzgm�>#"PwCn�=�|r���d���x�8�䳸K�A�=�oXVȊTn.R�(��~�lՙUd�/-��mYl:&Rlҙ�(=�*4H�#Q<�w��J�փVj�7�EQz��%$u=���]���Tn�U��Ў��������Z0���b��[[qLW��b���vB�<0�^��tUx��GX��������4T�@fm�%�)����ׯ7�z]����^}4Z`7�D�q"ı�;���@�q�E�2�p~\?cz3Y���w &��0vJ����EZ�Jy2?����6�}��K�F����Z]K����ʛ��638#�l��/ij7�c�כ�(��
'��V��q��G��t�m�̨���?����b��$Y��9>(�,k�����}>J�e01�/��w�V��3�֧Wߧ���-��;uɖd(�2�I!�N
{;Vq��%i::_#�⸲x�{���~�z]@
^�B��l���� VOB�nm�����l�ş�)�u�W>KG�
��)䭪����n-⤭>���
�B�~�
��#�B��E��A�������cXK����S��Myt�:I���*��|;�Ⱦ�~�P��5o�=3�_�<14���X�j�N�n�fӐ�8[ t�L���_r�3��b\
c�Vb-Z	�1'Q��J�x�d닕�־ZR)��C�u:H��/8 ��2x�Q�5w[�t3O;j���Lc۪�C�3�k��VW�+��C��X���ӂ�����G��F�͊n�O �[�q5��w㽉�%,D�س;�0�"D���S���ovt?�3��şj�e\��_�D�i�Z�#��e�����~��bR�k);�������{ G�!"ͥ��ovQ
h������Y6�	I�{�T��w"(�}ޑ�
I�b��a�[[`��@�����8�|�z�l���>A��XoԌd6'$��R��gx�bNp���[�q�Nh��<��A#��3�,��=��u�^t�yFY��40�S��Sq�렌��E&>�Ĥoԍjiűa"��'���Y�#�^^���uY����0������6�l�%or���y<�!�ln�n�,�gW+�m�n&Y~N�R�b*ێ��|�ہ+�<U��N;��)X!i!���_��Y� �$��&���.J~��n�+���]�ܿ1�cNx9+�D	܉�T���O�8������_��c��b�=����s�9��G1�����֣��JO�����3Z�P}'��Z�S}��cr��䁉�/l�o����t����Α+�mY�R����٧�����,��[�SG��+�R��[y�� l^��.uvypm]�x�A����{�?:���l"@~gI~ga����n�o�p=���*m˸��L*�������B�Y	\A<����8��"��^���\�0�_�8������I<�n��|'�I~k�L?�VQtron�1bK?GzX+��r��ÇP���^�!�ԝg��[��7���C��Ҷh%�ytE��te��qU��v]bRX�d��kv.���y�ܲ�s��cW�E?�</��!����ӊ�;�4G����u��nѼ��͆2��E�5y�N��ݪ��T��]���U5�����<9�CO��I�SYd8��^1��G;b<��zfk�fk��7���fY����F��g��r�zK��愓���+��'�.��,���,����Id����uu������D�(�B*���~FcF5[�h�-aΦHіԔx)���(NS��;�q�D �CS�aY�����;�esVO��L�`a��,�-ϝ;��2�a���a��i�ˆ�Mdӎ1���T��TL�O������9�9<��S�ɒ�降��q(��7������VZ�b��.�����y�= ��-�����bG��Q�6J��F�����L�=���R������X]���#1
5�z36܍���U�ny0�,��Ef� �����P8e6����,z���!A�+j�o>�e��C����B�̚�g��|�@m���^��������xL5ή��A2KN%�G�����d��EE����`�6�Ʈ��ў����z���E��%"�����:	̿�aeBE���E��X��S�b��:����EǱx?z9��P�O�E>�ϩBNƺy(mKN�l�#у����><�w
P�fU����,��[��77��ѯ�${u��)zM�F���Λ�e����U��G֞��=y��'qm�G��j�1|��ݠJ)ʃw��=�[AW���A��TU夂���[�.�eơ�}�zJ9�+mQN�Y�U�ם.e��O&G��ŭ�Q�4Yxܩ���L�V�K1)������I�����,��'8VF/2�!I�z�Y�����;L��`�L)b�D�w!�pH!'?u��'w�ɕ��-ɯ�yI���q�b����W�C�~��6�I���e5��z1��֕gq>���Ք�:�d$�7S��}s��2b��u�F�p=J���md{�LA �`7ZI�<(��� �H(z�E��j�����[dWQ�ѣ��$`�0NS)@��Z��`�ԕ�u{�6|.�ol�LI��JM"��-]�_�m�'����	���n[d `@8-�*����-���`ƶ6�pf��"`0�������?�7��є�sQ!y�+��KeOi�lr4��cX�3#���Kfs�j�tė��ڃ���z���&pO�r%�}�.���󐎽o"��<<P!qJx���[z�RS�^�U.f�'</f�oq�56Gu���\�R�nvN���_�7��a�q�������\��b�ݳ��L^9���ᩇ��~x���!�W�ttI\��?�z��6��/tO��TM�;���G�6�Y�ҳ�9
��D��O�����@��_	39�����%���%��7	V�?�_ �?��$����T�'�bމ@���%��7V��̂��(��������@��������+t}�IHHD��:�}�������:��0���:dc� ^����A[�g{C�+�n�T�����5�L8��r^m��*��.�DcV�OL/�K?'�z�l�?�3�yl�������5�����ݠ}����t����x��H�[+�*B�bT��ߑ�_t��N
	B\Sh��g)"�)����Z>Wd�4f���>�m�j����318zd'B�%��ܞ���W��-�vE�^�m����)���ĵ�L,�Z�30�W���U����[7����������P����е?E�Q�\q�_�ɑ#�j4�W 3��@����ϴ����9�Uֆc9e� ��;ۄO��c��v}�����Q���o���,kY�M>	?��`%;��y
P?��gg��x���(���7gnK7�t!�� l��J�=˔�VM׉�6�^�M�ߤcd�7���=�7����|GHdJf�p4)p���]�* �y'�V�'i������URQǎ+�U(�Wg���A[������9�}��y�v�c��g/��!����o>�m��㧍�$�k�kM�'n�m+l`&�E�=�e���o�1a�hi�
;��,��K�m�߷��+�ݤ-�P�_Q�\���W�AX�.������H46�x �{G�6�#����l��\��kS�~�[�� �m�q4�%��+��$����,ƙ�[�+�WW�=���g�-�r��A{�W�W��_ �24��ĹW:�����}�&赯�݊o�f��u�{����0��j�l���c�V�m�v�����ـ�7�e��B{{{�~����#(�l�o9x����ݰ����{FK����j_�҉�f�s���j�V!�J�wre��reӗt��f��3t���D|L���4����/�
��V���mJp GPh�� �y�����b���G�����cM�i�=� ,�`υ�F�hj"�B��?�V�ޮ�H��Č����Ə�)q�.��p�.�S?a~m_�S��\2���lZ".�/��=~�͗����9!�n��8œ��u��1ѯ��M,.�G���l�Udm�?��{�����oj���Ɔ�0aV��]aV�V��g�)�s#/1t��DG�yQ���`���F���Ƃ�y�� �֯�+�W�j��r>���@D�R�2���c�j�{�x��V��/�4T�bu��6l�JT�8��Bx�D<�F����1237?�^	���;�>��z`>�j�	�δY�4����5�m!Ci1��F�yЇ��V{�����6����p"�c/e}I����n�G��bݏ�V���z[ܯ�'�9l��7G��:r@�6�|���̇���\�&.�k�Q!_���rsm���؞VFdwyQ�lA'�qK��*�cam4�p2a����G��6���'M�ϙ���?:D�*n��g���ŗ��Ro��X_^
����xnO��Z�-"S��#��׬�r�zT���X�d�$�x�}�����KoS�,dm�����D�x��t�┬����D���1�7YK��GP�V ;�����vu�8v���$W�4b�� ���D�|�ul ��JN��4�͝�%��Vs��p�n���mZ��7I��ˀ��.�&̺��W���m��H�X���J\c9�0vH�MM���r����\���1ă��&�ܢ���ty,T}����ܥy�CWt�M�l{{�z0�zp¤!��u��CĤ�X>��b�`n<=�AB�ki�5}6�=u~�V�7�"�t�m�p����[���=e����&og�V��/�p�ז�3b��(��X�E�e�6�Jǔh��m|.hXr:U�HPml^�"n�B��I����X�`��N&6���,��_�޴�A����a�4r�.4�/���>��%�����L�|��5#ٺԶ��oG�d�EM��U{��������=&�?�y����/C1�ĿԶl�X��FY-�?��ŞjD���J.�=��g!��i4p�q�%堪�\�k�]b�#C�_��t鷓�>���*q'{����%#��^�j�p�ޞH	<z�/�8.����l9�'_�Q5��Q2l~ظ�ͰMS�Q����u�������F��C�6�������܇U� a=��O��͖Pf=fդY�>}?+C|�p��X��Y|�x����7bw�ׯw��K�.1���'�vUt�I��bTcUA���(�Bv�,��3Y]b���>Ԍ�x��Q���v]�a_}�q�p����U{��q|�ك��ǸMu.we�/�浜72̵��2k�'�&,y���v4��Z7De*�����b㔸�Ƹ%;lBq�P��ٵ�N#�O1K]/��vA<�)`<���G�L�8g
`oQ�:�?�p~�Qcx������Rx��M�cڪ��~��u2�y�O�|؝;� ���wF�u��<]�������s�7V2���a`e��U LL,6۸#��S�SSSV}��+�Y@���{p����ߛ
"u
��R����_��qȼ�^y3Qh��
�HNE'�w�þa��x7�R�B+%�bu1)��O8������b6��۞[�0��z)u�bOO����gb��HM�o�;����U4^%���8l0ף�g?��x�:��1K-�|{r�e)	�+op=n,	�yV�(�*�֍��Y�r���sz��7��Y��A�57����>�o�D�aм������֙Z^�%l�Ͻ!����t@J/�5s�R��݉]Qy�f!�j��)����G��楀�P�v��AT�c����]F�����*K�V[ .*�դ���'�k��b�~Rғ�Vpb�ˇ��kMV��4���ҿ`��WM��W���Ɵg�k*�]�=��43S�t��!�<f"�K�ؿB�V�7�X����o��6��Z������=D|�:d�%�_ߥ�Bm<c_p����ۚw܁@��3�@��~�ǟ�5��.I���$ޤ�D��R{����r	zx��J�z~���y�nLtKWjZ�Iu�2�G엣��,�E�1@:W�2�e�B�� �TZ���p}�t���I��;gk.��Z'�w��\tqG6�n>4������Y قș������#�1�~|:O�i: �U�c�A�!\���M���.sO��f�}q�&*v�� ���/�5Im��Ffl}�ٚ�_To��ӼR���'������\J�Y76��~�<��m}XʥC{5  ����mԤ�+����]�]�Ƶh�H2W���Pf&�I�g'a���"������-n���M�R��`� {����8�����Y@�Q�O�w.��x�$����7��ЉcK�S���	"�n�_g9C�F,���Aπ��G���0�'K�V���sA]���Pg!���4NG�>5q�L]��H��}�w+��>.Ԭ����xB���^�BW�U� J�U���h �ۆ~GI���8Z��P8�m�ץ�)E��G�ڞ5M�א���ęC�K/t_����Ԡ[��Nj�*�w[�aI^~�@��e�h�=�NMݲ�=�b�JϽ L�Q�3]�$d ����E�v���"��#���R׫�7�Dj� E"�������u)��Bw���Љ9ð1!�;�?��4to�a�����X��	H��]�փ>�µ�50�"�}��E.]9D�&��1Us��n�jІ�D�Xm��7��بǷ��[��7)M���D�Yl�.J?�a�q�ٯ�]H�����J�SV|������	sUe�(w�&N�^��j��1�g����ɪ|�wƛW�7g���i��1>�]��C���O:ޣ�R��*��P;�=&m�rn���0���w�p��#Zi`��.�ׂ�W��S�*�6���u��y2����ET����Ε�5DU�k�.�>��NdAI���wΉ���Q|�`�z������V>��1������M�Xlg�.��F���5#�X�N�H���ȓ��3�d�#�4�16�t�����n��U�����!��S˯Z��P���n
��(�+�߉��f�:�f5�\I���>d�*�Ib���Nׄ�����SY�TA~����0����̢f�l��NH�ӧ���v��H�q���TZ�w(�?�E�o�O,��tXo�ay"��aL"�?���9���!LO.Ht��Y&�|����M}W��p��T>�m{-e��ǥW�Dͯ����:镅C�����x0?���jML&J.7���cU����%���3�i���$_{�M3�M.���ۋ�|q��� MQS���M��x�k1������"ቡ�5~�G@���?8�JCB���6����%�.��A<��$Kh�^���y�ܼ�/��{���~���Cr6���v�w#�q����^瓜:K���]Ľ��	�����qM�sE<�u�?�j�Y�h��E�̷�n��%5�p�YnE^[n��3�����ƺC���O�!��-N������譡��a�f�"w��L�ݥ��,f���a�.����i"�-����l�������EK�ʃH��;u����N>}�F�B� ���jHX~���=y>�n>V���{ay���l,bMϢ�_���7dt��x��26ͧ^0pS 6��5�w:�g�c�(��kn��6)�x���3FFN�F濧����~�����"+�� ��]������e$�k���?��&�1����5Ɵ�:�7�*2����p_��QS���/h����Q��>U�b)�6ݶi�:�4��h��S�Rҕ`����бe���R�	�c6ӏ�z�o��gy���%��R^�+�А���♅�]��Į�.:3*l�H�ם���4��·�|>T���T�+QL]F���q<_}8EV;�]�b+0>ouqq/d+$6~�, �)�`I�@^��޳|�*l��v��d�`_��@\�sl�����WjeR�.���{I�(�%��V��N�BvB�̜c���C�v6���W�y8�C�?���#4����QO���2s)����k>c��Nԣ�%R��;���s���|o�֣��Ӆ�|5���gG!�������^%��*l�S^dɟIg�u���O�G՛#tN�.z��M��8���5��i����ό���y�ȥ�U��,>̀P�7�Ɵ$�[��n�
�0�*OM�5��r��ta���7�rZ��@W� ��Kw�z�DU�g�&�'���v5�Kd�E&= �! �dk��+]a��⏲�W�녇�t4�~���+�3��j�Vr��9�LC���Q�	)t��L����(K��T�w��/�Ԇl:͍sfҹe��E�WK{�BB7����*-���e&��'MԱO�ؚ��x�B��鉲��"�K�k������MK.=��p1���y�=����PH|hr�b,^��Ϲ�w��l�b�f6�<z�Oʽ��қB��$�Df�7�p/�|��s�;U�1���7h^��V4��?K㈿�������N�D�{��)�����_�5���o-_#O��SÕD�c�~hg�䢸�O���J��>��`���|z�� ,G6�iɵ����pa!,���P�LOJU6�������j��!�����&�,Dw�`�N�YE��W���w	�d���'j7oa���0A.�coKl�����b��[^qtc�k�@��LM��'�o���P��	�;���Gl:`����(I�e@)(O�]iB �q�W�>���K%�*�6t�~]��k�ub� ��;�����N|:�침��{�oU����'<q�$�T>�����ys��N�R
!}4��-t���Ѵ�
h�?�e6g��Z���ӫ�g1[���.B�B1��3|UFf#Dڋ�by<�K��B�?�W���3����d�M�����3a�	~�o�!w xh;�na��Ĵ��A�Q���)%�#W�`&Uǿn&�D��������MvN�R�U���G���Ն{��9!!K3�Wϟ��8�~̲{B^`}���j�k�d��>��R��?���y��Y%>Xq���pGy�j��I'S��Cg�*��D�k��=ZP7���L��\�^m��p��UH�%>D����$�������<~���#t,��U������M�	�$�B%�7L�p�5�����J_=pz�� 0����/��iĊ�W�v^R���,�nt+�A�Y����-�%��g���-�x��vt4z����[�~�����Z٘���2 E�*ݴ���o����L3�M�*J�և�ɠ��R�8�9Z���� ����Ak�����P_{Io�^	>�v�p'X�����������]n���m�L]�̤Ȭ�!�(SfJ����1��2���)���2Oq8���1��]�v?���=���Z��z=_�����k�j:\Tأ^/v����uE����R� }G^+il��>ɀ-,��su�nl���R�ŏO;+�[��[ ��D4�������s�8z{-8賡a�/�>���~
x��$?�7
NF�rg�m�B6�=�iz���Ʃ�����眵�KtZ
���:E����O5=�dm'(p]*�H���B����ss�V��E�9��>H�A�H_x���I�s�}�m�Sfqc6��/o����C�p���J�u�����=���/8[�_��-���P`>�iKp���ε"�y���`6!���e|J{z�ʂ��p�ιy~a /!]���7�[�c"e�/6���(���?����Ǩļ$��-��+2DL�u3P�
ޡ�/Q���z@Cu�V�iH��8�P�{X$Tۮ��?uj��^ps��[WDO^*��nN����%��C�gdt�g"��/��xC��E��%��B��S����ŵ�z$C�b����0eu�9��\t<����5�=g2���+�5�/��3��e�9['a5�G9���7�뀩��.ǧ �O��]2�هac���8h<��8��腂-{���.�=6%r�oo*��"�2;�C���E�J���Yl��6
K&�;`�=���f�4�9kE�=��}��>�rO���}�<���	�R�{AD��e%�H\fy"��ۄw�f�i
�E�梔�tv=���~����}�zd�^�i��}<d�5��kg��Q��j�=�{�P���0�6�1��lW� ����BH�3�����f�Z�>���s�%��\	�Ǖ�LOd��ٞ���p�{J|ieI���5p��Ԋג�UU"�:F#�n��쑛��[?��'� X�**�p�O잷m�z�lA�k5�D/
T�/J$�+(�P�J��Zy��'_v�fХg
�cQp�^챙"�^{]��4Z{IDi�t�{�^����uD�v;����K he��B��k�(3��O���}�Xk�[�wZ0�(���[N���t��9����4?WT�x�7��E3��)�tW�_^�$-~/�����U@;B8�����ʵيhx܊����,�kU�������mω��, g~��lf��"Ҹw ���,l�QT
�$z�~��r�.$P^ ����߼��U�C��\��ֿe�0ف��?��d:���&�m�`2hǯ`*�⬿oL�!ꣲ�u����R�ZC�ݲU�v��Ր���@�\b8c�
��F�}�� �2�q"� `gO���$�y�#��y�=����q����:�8g�`�t�.t��B
Ȋ��S��4}�F1���6����HK�ٽ(W��W��c�)����n\�iȗq۬��ת���.�x��g(7���?./=o���b��)�y���R�bL�	�ѡn�۟���kfC�~�'��S#��p+Ng��Õ}���z�I9��?��^��U�2�m���1P���=Z�a�l�	�:��>�Qt_�G����P_��[�Z:��ON���qe��G�p�^ n���\�9R�]Gmi�V�ȯ.+�ߡ�������V��
@ș�w~񫋂�5�����{�G3���c���{���V��/WdB���wVQ����"�h ǭ[Ğ�zY���(�u8S">E(n[fɷ���Gr���B���aZ)H�N+6r�R:"�e�F� �W	u�Q����S�6�V_H�?j�|��{V-(N����(��:�|�\w0��Z}]ۺ�{����#�a��ur���z�	��W��4�7�)�4��B� \j�Wj��7^������J�θ�<�7���x���p���V�>���.?��u�
G�2놧��!��;��C���+�ƕt�3ٝ]���
ؒMk�3�_�M����)pq���Z��E�U�{	ɑ����Ķ)����dm5��h�-Lz_L��b�(���/N+��+f؂V<J����t��u��@/9j�DWg�����%&��D4�w���V����t�1�l����A�ج]���S� C��)���(�bUT0:�?�
@[��+�8���e��3uG��u�6t=�_���N@��^?V2�PI/!�v��0hX���솘��<��>gJ$��h�����eFھ�%!�G�&��R��/嬝�C��O��4/|G#m����i�&�f�D��^o�=�A��ske�c9�Iolǣx���{jq�=���9o��\�����'�,l|%��� �[�@��$y�������L��E[c�L	�;W{Z1䱃H���3DM��i4��1(�G�bhf��
��x��x�� \'s� ���G��Y�D�H5����G���Wq��#���"�#їP_�d����7� �d��X��:�~t���p���E\�ФsxFF}th�$8���7��7�e��:�Yw�� ������f`�&	�˷;`o2OF��X��� -��8�}�$)���O*�H@��HM�Ϙ�J��Ģ�w ��:[f��E�����^�HU�z��0����9B1�S�T�#LLv�{�U�lRT�#$�(7}�u+���C��N�Խ��B�b0]��JC~�M�C޺��t���Ǫ�[�#㵊��ď�3�(����S�ſ��eS`F�hҹ"����e�Ѽp������(
���	W�*1��v�`�gR�X�������?��� z���gT���L?֘��T��m��B۞��v���9G��]읠�5dzFd���`�������͚@[QB�g������A���M�a�#��"!�P@���ܜI��dQ\x�F��.�f�dC�J��P����]��
�m�����������;�.���iq�yQf���15@5[c�rqT�hх˙��J��c���t]����M��w��>���\�-� ����~��n���`���E\�*S *^�6��-���:u�L'X$)�ג����}�K�q�;/���/�
��"<�yzgBbz{�=S�E��itz�[���V1�r�U�2�7�1��:�΋`�P��b9;��[��Q�<�Z^��9M�vu\]�:���W2�]5U�i����t�������	�؃P���)<��`ke�m yF�K�s �_�멿�\�c�t�n����)��vE��??��`�ǵ���ygi<^M����;�~7��)�%���9&��MpI��,ՃH0���gw�:����'��ǟ��S5,���sTM'�61�-D���q��Rcop��kQ�
FwzT0=!�v:'y{$����Դ��w�=��V��ơE�����^����_��U�c�*e�m	-ά��D����m�TI�cO�����n�	ܿ|�ǂ�b��q��s���l�ڴ�Z��q_��EH�.O&����v���w�4��7Z
f��D�l�#/���}N�ٮ�U�:����=9���-H� ��V&��_L�l74�����d;� ן�+\�5�9�]�¢��\�b��F�\�-U�1w�	��aDlʚ[��Ƿ|d*��i�����V�8��\'���y39~�@#�'fz�a��@� �aH��J��M���7��M2{���-\��70�����=������,�3I��nR7�I,�,zn|
�Pe�����/��:��ͧ{�VzI[Qwn�jG�Ʌ ����J]�"]��T���I��7�+<��(1D��\�D+�NG4�L�%^�o0U:�����P�������E���3�otB���@�9� �B(��жD?U��õ��`�gD��o#�d����0v\21����s�d3�����X+�QI;k8Bޜ&����ǳ����e��y�����Ƙ���vXl����E9���6�����va��7�=��2�Bv��Tߺ���/k��\(�����%�6)�u&���{{cv޿�P��x�o�_�(I��r��??Pz�[Nse��a���^��7��3|N�<� �g���!Iey�j��w�B�'Bb����ph��+�Nx@2�����,T����f`�����â�\��|8��JKi��n5qä���i���UT�CEa��4�]"lP��K��V��&S���r�����AY���7��I���	�1��)�|
K�����3�an�>��2��h�3���#�'!^��U���ij(��E��;�Laz�"ӳ��BQ�]���A�)5�L�s��T�Ls1	����m�%˘�N#����g����4~���(+8_t�V�\:uL�|2>�=�3��	ix��K���qm̔آK��;8)r��3�ͽ�M�~�\�'xF�̤E��A�+7�L��kU��sʠ�V�ߎ���{ul_,�]q 7�\�E�hZ�T^f߮���ʩ&��E�^�,�ߴ���S�f�ה�������>$�n���qgS�l�-��g����N|�}Șk߶�V�DsE�����*Ԫ���?2/�;��K��U��\jy��'U3��/o�o������:�&��R�\�RK���Mö�k�8�v����H�� ?T(rf����wiwU���[�TF�И&�9U����	*�����d�Qg�DXP���h�����DC͚���:te����3�ߓ���:v���󫮮�l�ט���:ԕ��u���8-�qӦ��@�4].��f|NĦ�*s8��Iz����:F��xDԔ�6���hb�$��5�9�P��b<e.�@��E�[uf4�*0
���s���i�(d|�w)�M�dwM2���W@)���?�#�e�ܭ��[�)6j���ޑ��a�rc��O�[uf������K�D޲ �e�}�ũwʫY�����!w.��teb�_mX�� Mb���W4�5�9"��֝gl]iۑ� ���A�)�^>G��Z��T6`� �zz���k��xv���Y�(�I<��d�fd�P6P�Qk�2/�y7%����:�:]��Q���ȹ��R_Q>�z�Ӱ�N�~�wJ��s�ߍwDT�6h[\���I��ҹɎ�r���m�ŖE���v���;�T)�X]S�]���vc����#6Jr��dȼ`u���G�j�gq�	�s�|�C���.ՓB��NS�EYt�IQ��!���K����q�(��W�s���I����7�j�7����������t���	�^���7��Ê��}�pG���)�X,w�$�����r�^Lt�pd��\�����ƙ��9$����̩�+�U����j�UD�x�0d��XU��g8Ը�0�����[ID�PL;�_G�#E��sS�bь�A����X����Sv� ]�����v~����wV1ErHk^���n����đyCMowJ7ݠdr�I���Y��§��Fwg�W$�jU�=��dJ��{C�4���}NQ�'�����i��ɚ�}�7����A�3K3p���e�L��c�_��z�0��UDG�ot�R�+q�f��$�~�T�����^0֒��g�A����rs�m��߱��w�����3{�
,n����P�"��L�l����>��t
qW���w�,Q��K"���Esi�h0�	EKE��p���韓��z
T��7��g�ly&Ip0v�_��Z�Q�jqn�7/± �9;����܆�O�[��K��&RHA%�wy�1���l�}�O0k_��'΋-���uE(��T����H3h�|�1#���ct�|˹N=&xփ\R4(�=��1�1@�())�P�gn���մY��0²��cPl�Fz�Q�v��}�fp���3�jȷ�+���7��l��f:N>ʭ�-#�HK٨[����?��a �WO�U�^���-~��w4	,[��&�>� .�P
㩅���L�����嶫T�T0��*K e}V[���"a�5;KjP��d FW���㒊����ʊ�Y�}� {�㻼$��(n�lw���%��C��c�ؠ\��p�h[^I욹HA�����R@�G���3��Ӏ�$�����okdP_x������ۊ�	�uF����ϩH��X�(���3.��sUvQvxq5K ?1Q�+�{I*����Gs���ec1��74���.�������^�MB��A��1�G���RI���ސ�َ݂�J$a�ݸ}C��~iT�͙��u_�Aش�hʆ��>XpndxRu2}��0�Z:��y�����L���Bx����z��*������#Ώ�F� fB��N����_����R�S[��J�DP�+�C�|c�!}wBz�']�zPV~_���K�:�AeX����*��}���?�+OIQ��=p*��
���Ƃ�f�B;P�k�����ϝ�����Ef�~e!��e���7
�������:���I���=*?5��ͻ��t'�#4���B
�go�l�>/*	G;���,y*�����ցf�7�[�� ��j=J�%V�b�=��ѧ�J�v3��1�7܀37H�Y���ɱ|���**8%%e���|9�[3PBd�spi�N������p�|@^cb���4&�36����Ow��磑V�&��4_T�L-���w��|u��&��~�h��^���UZz@�~'\,Ze�7/�^: �"!w���ja��ĲE��'^�����Ra�h��d�qʫ�1=�S��B*;9w&>����-�7�x������=xAv�l�3�_�א��:ǻ��X[��P�%LYǃ������r��Ie�������=��VlA��2���K����Q�M7����0�DWg��<��Qc��S�!�Y�߲��I�Y2���h+g�6�����E"���}�|Co]���"\l���l�5�����*�8A��gM�1����2G���_M�lp/�_�F��`�;�uU���~3�V%?��� ��dJ��6���c�N��n�ڜǣP�>��_��CD�n��-e^�tʹɠ�h���dĝ��גܖ>�#W��6����M�����FQ���_�ꮕ�M
�?|���� ����T�u��=s���|`�چ��V��v�������3�p2��W���V�$�Uy�E{�����l:�<��*Ɛ���(�A.~��WB��A�5j}ghY�~�1.���+�T_L��Z�l�O��خ�<��|�*BW݉�ο6e�8+-	R9pXy=�0��:������b�.[�OJ�脤zc��6����G���qB]�UNf�o��M���Ԑ�;6M������y!����$Ѝ�`�)%��5�a�?�:t���1�ѣ�I�q�#3�?�H�j�Ϫ����j�9���������ysq�5����aD\$��#��ɕh�V�.t�'�Y~�;R���S����c��T�r�P��{]s��������٧>"�?��|��v�ˡU+���n�Cԕ''���8ɁS�3A '�����d�c�P�A�s*���sm4U�V��K#��N������%w��:)L0F�oа4���F�Z��
P���L�U�M��s��ѓ#�O(�g26�6]&N0��I��5���?�!��6'?�nQ-�:,D���+��L_�X��VS��_���C�5E �؅B
��6�a�	�M7�McY7ak�Y�P���X�mˉ��K���%2vë��Нxi�0ߠ�|*_��(W�b�nm֦T�)�7�_Z��W"���x�D߁�,{=�H��?W|V�e��.'�=��y������YtuM\���/��r��Z�E�!�у��>�h�[�5��j3o�:ڋR�O"�l�uoZ���7��g&�rq¸!��|������Y�m����z��������omN7{Sk�r/�*T�r~�*+�J��?�~CW��������P�ʲo�Jw6�ɡԭGrzU�OH���/�M�h8����wL^�������V�^W��=�i�Q�g�q�7����h�՘EI���_��FN�L�^v}�J� ��%t ��a�aY�%-򦶬~��d4C�����x��5o��2Mϛ��Gf|V�M��������+�Z}|�}�����h���>��@��^�C���j���H/a�����<�#��S����m"S�)L�T��3�2O���A��;����rUUmЇ�*�F�/&�P��)TU��<n+:,���>�����Hj�1l��*>p�ĄD��ۚl=�q��2��K�-�y�E0���R�i�Hg ��>՞b�Y�ﶫ���iv��՝��\ѿ΄�Za��,#l >tt�g�̓�zXm�^����f�O����`O��z��A�R_o*�")Q��K��_VD`7�wO�����⎴��j����r�7|�Te��Ff�$�{�7E�X��s��I��ZuKҿ���Ę�.vb��T����:s���#W5[��ݔe�g�81�s������K�K�_�\�%$/jH�O��nΙf.��v�U+�N�����k_�,�]������U�k��/�c|VS|V}}��.�{v�rn�蚬zJ�f��5��԰��";�_	Z�>�H���n�b�<�;|*NӲ��1���@��L�RA�e�a���EjY6V	V�/:�G��*�"g�N���[�W����od��7�:���MI^`q��ԗo@��։M�5
km����2��0P̺
@�IZ0̶���>��l5A�U6����f�<g�8��t����M3s��ZԢ��6%ډ���ʜ���ֶf�����h-ee��/1���_K�vF�8�g����qڝY�p'�zWI5@� zR��eM�K>�T��P��t\��n�sz����%ܿ6����c���i���fO��q�������Ykn<I��@]��m���O�5u��A��Nrb�9��o�e�\t�Zm�x��u��Q!P��][bӃ��ٽ�\��2C��K��J�2;�./�	�f��+�,/[e�,[u���5k?�
��s�}6v$�|*�q��8��^jz�:��=��2���s���k���~�e_���yp�ҷ:��|�tb>�q'@?�NPp��-������T��h�	�g��K���y^P�D2F�}@p-�jOK��Fv������e��g�-]\U`��F��D8�<�1���z��v���u�̢hw^��M�B���:�i��y�-~/,B� ����L��Xޣ�~oc&:����q�s?ێ�q�h�8[ad�"�Cp
D#��x���d�H9�ʮ{�>W2�5���i���^��|
�/�
ְ8=��Kt�v�:rd߆O0|������W�:��#�AC� �tqG׿Q��g-"'[�����긵o�)����:y��S������ ��ܯ��������兼2��m�u�&B��D�$փ2F����!N&�qA����#�K�G����?V�j:���
�:��I�w�����Ȭ�b]0��>��M��??�̥����1��������R���c0ు���m�?����M8�8�ghlE�_�Ə�� AO��z��h�A���O���S�l�H�\��r���4�Cj�B�8�N�с�d\i��4��駔��&�RPo/e��t�XJH��Z,.��8�ԸË���SD7$v�L���X~&�8[N���s̛�#��s��p"�����8���<�FDD��Aj����g˼�saJ[_>�\8�Dj�Ճ�?~������������J$
���NV��w�?���*�(�äƛ7��;(p�?�'����]��W��]�4����U�p�Pp���^�^����ܿt����m]].�C��H�Qؚ��S�;���FH��.!�cpP�Р|)���t�
�gg�$]��K�Ŏ@�H�s@qʡ8�`	YW����5D���۝��ѕ��Α����B��N��O%��N.�445Uon�Ʋ�Щ�$4�������ǅv_��+.C�T�zA)6<��uu�5�ޢ��fU�]$��􋋋ٰ?SCH�� �+��P�/��W�9`��LS~!]���	P"p����k��-#=D�nz��ťW��5��� \܄�.�@6I�1��Z}�����Hc�2{2�WZW3��& � 1P	1J|�j�C�u[�;��@����]3�}��@��M`��o��ӝ�3M�D�C0�Ll��B�|����a��e3`��P�+�d�I��F�9����Sky�h�_�VG�J�b@�6���P|�0�Q9|�:a��]xZ�@H���}�7H���cmm�,BY=1�}o�9��ty�H$�;w���{+dI�Gi��m]������5��+���p^H��e��2b��쬬?DIm��-�t�=,j�f�J`6Ε�iݓ��b���\m����)+�����G�¿a�x��/��vBӄ�B��TPXHOj�V��=��ÇH)6���M����+ߺ�{��Sg�X*2��c:���jj��K�yS��Ǐ��_�jY���j1l�B4��n��ul�^�����4:������G
����}а��|�m�+?�]�?0���XtJ���3R���+��Gܿ)�hhj�K��(��3�3m�=@0i�jbb�+�A�O=Gy`�
�!��Qb\|�bG������O�<����
I�3}��
�"w�<�G�m�:l��>^��T��펙�|���&W��ɾXۏA[2��h4��RM�3^��\b�M�W��8�}����	��[�����<�Y/)$o0	��p�S�2�pLj(@F��$�l��Ҧ:v,���6��klj
��ӛoc����q�%C����BA�*���~On]x��YZ�~�f��i{���^�vs� ���h�&T�0�����w�=|��C�Q�iM�W��?2}�O2W�X^�G���������R?@�W�Y~5���Zd�PAMԑ���9�}?�h-�}cEk`������BC\{�Y���֩n]�A� ujr��Y�,oƴy�aIMZ�k
�Tq,{�P�	�+~+нl���l�(�����l�9��I��|$�w�@r9��m�_'�ꨧ3YW��<J���+����=]�}}��F���~�����a��	�\8z&&�ngN�N�)P3힚-���*�����ع����8�-�F-�빜Ej��6w�nі%�.
q^ӽ��������:����T �8f	�
[n�+���(���d<��m���K�����-�{X3f�82����T�[W��\�|��5�t��3�6���D5�_Yzz�������h�*�-5�8Ja��t%))I��Iz�W��o�ځ��{����S`d�>N�(U+M.��~|��U��Dr75y�P��!w�=G3�>6��Dl����}�cg$ �o;Ȭ�o}9[U�ƍ�-�#-��$�Mhp��:4�e{�	:7��'�(?��܄��%�E͊ڏ?��2�p�բ�<�9ML����F��^6��c"}|���RS^ZX�j��~A�b���J#F���l�qUS�O�mll4p~����� ua͕��s7��m���%����q�HY���3�ֿt瘛8����+X�>U��E״����g�j�A[��]䞣�[����y��`��V��H�C�i��A��#,F���z��W�,J�F�����Ề��:k��7n�8WfY�]�6}e{444t�������ޮ�q�aS�� �N/��.����ȷ�n��6��{l���3R�x�,h��u�P�Y����4��M�g��w���˿+��q��G"�^I����٘��c�^�)��f���A���P�R�hS�8��Ӈ�
�|1�ف�����1i�ò	6���=�Q��{�p�&���T���� +���F���l�L[��q��=w�v����ʰ֘�^^>�j8�=sʚ楯�oW�����~��`7���P���p.j�IF�(�<�z:�f��?TU�2^��K'+��<���e��Aq�����ZXI����{�(�~��_M���o��q�t�W"R�д�G��r���P�.)}� O���j	8��gce�WP0�X]Sc��\D�uez�&DI���fH�F��ٗQQ�e��|׆�Qt��?�c��8P���C�jum�H_6;7׾�H�ҥ���rM��R��!8���W��H��(�����ӞNߎU��)��*����O�	dڨϧ98n�G�Ke�`��1����� |X�F�yHH@�Vm$y����9pBd�o�)(!���s�y�x4��zxH�ٞ�C�)����"�	l헮W�����8͕X�i��c�U�%���(��h�9=��]������	�y*�6S�|d&�����A��A.���WD���?)�}�?��\'*����=�:�-wnR��ǟ�J����$>�= �v`���A@�+�)b��X䈷�wɫ��
7//�G�<||��zy����if���x��M�%,I3�b%����ͬE>Y%���Z��/(C��pۚ2
J�q�BWl�n��&�:�>a�Ɍe�i��9�}���� �r@���
����gzŁ��LR�VV�|��:LWA�*�v/�j0�+���Nc����8�o���r�S����qP�ִ��e�"��և~}�p�ɩ0�$�)�� V%�*)�
�+b�DV�HRt��	�g
��&�؁|$� .�E<��
pi�(�D3O7���..&�N6�X��<m�z^��׍vUi&�U��Sˬ���AQ���r���l�`��Fڗ@�O�
��,g���l2����
��9�*�j�IM`W�+�w#+���{��L43U��w7*�%��V�dYq���� 0���Y���p�豞�)�i11q#H��3���[W�2ɓxPR��s����S�{j�n��j�Ν����1W���	�q�	b�п{E��{�;�i�$���t3��[��Fku�Ť
N��H���٨`�uܸko���>�9E�)���A&�I,-�`
�z���r�>(��2�Eث
����rF�XܗZcx2E�cʛ_Y�� �6��5U�QZ΢�
����Z�,�:��p���i�p�:��$�W�����H�u�LYm/��1�4��+fH��6QP ���2�\[��hXP:ʛr��[f�&i�-�����*��Gq��.i�B���(Y��O-6K�x��{v�F���j
��]��g�Μy����4�7xFd���?((<о��z�ʝ�Ov�8=2����Y<�s��q��@�4s2��6~�+0;�Ñ��}JO�"��:��@a϶�5���er�.+�qG����\����é
\�������"��G4R�t��ߺJU\��Q����";'�7��]!		Ɛ��#"�7D�O �O�c6n3T��b�kmW�þ����ʩ�X��n��nsq��A����{Dr�YUa, (H!Ow�>`u�^����w�d(wA� G�{��;�Z[[i�͒ѮI4�^=+��Z+-�{`�.�;o�B��+�azh_�h6��jO�CQ77�z���_(4�ū��;7g����� �T�t8e�<H�]@��q�Cũ�����fgg6�/J�,jkk�w��1��ǯQJӃ�4�D>�7��eh���%b��o�h�RK���t����"[��E�VZf�R��CUu��c:S���ty�]�e6L�U��R�jM��`ߊ��ȈM��/4�Ȗy��V�W���%|	�e�)+�	F�L���E��E1M����Sy��l9ŵ�+ֿ8��8�b�%`���O��4E����^��������0���� ��:���͕(�U�^�ZO�.eRv���p���T8��#eU�r�aאpK�\a�3x�S���,�)�;4���$�:�ye�����i�#���߹����HQv�u[���~�����=�<|\��g�c�E�P��,���R$�4g��V.l���1����G��F��{�O� >J'}��W A8<�L�z6�Zr#�Y]�_��s-�4׿���������֜�?��J%G���{P��E[ME (�Z�G�Ib��c�^ށ}�,
К���ͷ�B��\�Ə�r� �fcc���oS���ވB����eC��� ���*��4Ѫ��+ߵ�Le#;lq�6P��48�HhӁ��i� �cy������Cp���h:���7�(W��?J �1�;V��Yafd��(jQ:�e��x[N@�,�k?����s5ˍ�pC��i!�w  �Y��tog�(�I���>lS���&����l��
����V����2K{����C
�_�x�m�4777����<q��ի�S}���Ĩ=�O��:�)Ж^�>�_&��)6�RSTV��-9O��y�}���|)��h'��4;�w�@�v�[3&�&&q��8��Lh�u1��-��-����n5)4��𭷀+=�/�*
N�j���:�Jԕ�L�#����5�B�_���n���N%����Eח��th�o���YҦ5AmM5�d�\�{B�E�kK��90�9��B'�&���#u���ᗫ��Wb�j���B�Cň��R�C��SU�w�.�'�d��M��TWWGv&3���f1M��$%�,.�QPQ���#3��^�Z�����R2^W$���o�|AEIa¬�v>VEC�b1��q^]�Y$\;p����Oh]9]��m����6��f׸����e��8&u|��H�9ݛ���y'7�#UF1��Zb�P?���a�����=w�Azjs]�J�ͪ}�n��e�%:ZQV-����:ʜ�cQ$�a�]7٨f�X����!�ta�Gh��lfJ���;�cVf�{�.��
򱕯:N;�ִ��ǉ�`���Դ�J�AL�u�̄nkC2i��Hh�[w{��H� ��D<s���n�s���չ���w�ٿ�s�\F�ž|�`�@�q}4*6��k/̀ei#����!�K�0��`�h�v$%$6�>x���0�e�#˽nRB��^Ʒ��ȐI�"�i�8��@:w�e����\z�<ϻM�#�v�`��+�����ߡ\�s%�J�VT|^��Y���\YZZ�V����XU�\�qD��ɌW(5�Su�y��	��BC��|p��[>VC�x����N��:���:1QzH����Cޑ�bA)���ߗ�m���d�qN��#�:h�����=yi�#� *,b�qo�]�B���n�S���'�Ѕ������|J؆)C{�_Ft��� �8��ɺٹ��?w�9腾�a��`�%�Ӗ��o�Ҥ_�QW�ENW^��b�gPC�)t �i�~�H����x�X0rmm�#S��W�,�VP���@���S�"�,i�� �X��K�Q��8�n܈<�_G�.��l{��V��J�I���Ev����
��;m�o�x_)�\��B�e��_���3b���נ�Os4��?;{J_�r�!��N�7�_�X����j�D��;�T�rF3+#��*u�CHfj����eي0���y'�>j(��3���g(ՔG�x.����*QRTʑ�s����"�a��H���Z�(�-�G���lT��Z�wq-�U<�%���b�����/i�\ G��`�����>z7D�t�`%�E����w��O�}}�c@�j�?�ܗ��{�i�|g�'�UG�dRKT�{�+B̏�өl�B<��6����9��y������sǊ �k=�@�5�2C���b�d�����rٗ��)����S�퀌=�>NN���7�d0����/aAĝꩩ�rgL��(pg�;��%ќz}J7A����o��V�y+s�`��[��B���������Z��Q�J3�Y� KY���3_f�E~_k�N�uԄ��^�$�n�(��V1��8�� ,�2��bp�������w�y@��+J(�9�T2�gjb��ȩ�嚯���@�%z*V�}�H�q��C�HSP())�7�N�d8�
��}�@�b�T���P\(wgY'����Z}Lg����;���w|_�+������C�6;?�q�?j���P�q��[T�	���&Ȃ�Z][�<�U�C���;&��^a<uVP A�q� �u�;&��B���m�X!5ԹW���E�1��~�HGg��Gw	VL��~��Z���|^^�$�s�Wy�����`�)��e�^k�C��H�B@:�|G B�\���l��q:@�uj%�w�w�--e�3�:�\�1%�w�w��tO�2V�b�Nþ�'�b� -�g��x5�"�9`����*�z���tck��a��۲EZ����H�\~A�	�ls������L�� ��GHx���]RXDď4ekck[Q�x�laZ8::�h~)q��b�@��H=��� x&�,8�����1���$E<I;��S3MK����:5݌9��Z<���鮾����,.˓�<,�W>T�ih��7
	��V�s�_V6f�j�BxhCz�n�bj���h]���KNƒ���Fl���i[pmJ��p~M͜�EU==�
�)(�a��g 8�Z����"��EG-
���d�֘��N�
p�윜��ME�C�/F���2S����+���)��yצū�7�|����uH5�-��KIm�-��!�]����za}k��<��V1�S;��6��r��Ba|�.e���o߶U-fv8l�4K��</�_�P�) ����]���#d��hJJJ�H.hN+��ut|�uu-�V�E-��82u#l���jzzt�5<���M�Q��Y,��7l�or��XR����cu��ϊ��P�{�
 'LĿ�8A���VZ0By�t�j1����y��������ԗ؞h�'��{Z�B�O�W����"�ʥ��8:9��&�A�t'ڦ�_�VZT@;�&�O�S����q+q��3��Y&h�Bu�u��08`s�k=��e�^�ٿf$�r�!hU�7o����TVAlZ��⌄�	ق� ���jRqFd��)Q֘���������׬�uR��dJ�/X�"3�QI�Cn�6t"m
�H���� $��q�S�אs�R:�_hNPT�a��Q/9GV�)P��J����/����8�ֈ}�:iNCM�6�r�JM�{sT��m�v~~���	�):�}'�}VRS=F���F��A�$�Du)��HSs�8��� ���[�z������&�/��10gN. c�]�����1?"�)3K�(U^�Q@x$^K]%	K�KjF���H�8y��@���ylՙя�pE�CȎ�O�l��T#Yt!d�d�~|�7��4�R?:#�y��ǐ�,v���X�aY�Yǒخ�ޒ^{N(�1L�w/'�"�g�������"���o����I����ooo#����B'F� ~�UgQ���	{�"���,���vG�]���%�&f����RX�d7e�%/���i�Gδ
�O,���Ǩ�H�����>��6�V�a0�)P��L�˿X� .vgx�u�6ۜܟ���l�����?PK   bi�X��/F��  ��  /   images/24a65fc6-6c28-4ce3-80af-2bdea9058a0a.png ;@Ŀ�PNG

   IHDR   �  w   `�3�   	pHYs  �  ��+  �RIDATx��}��U����קd2)$@� �����T\�����b�����E,��P�� ���R$"���H�(� 	I������=��޼d2d&�̲^>a޼y����{�=�{α�o�oc�o����7������a�mlpL�X�h�2{���;��C����vuwT������M_r�G.3#�7���{r����S�ryJ:��l6���^:���4	�V%�;���+����_��W:�݇�xo��<^�̬Y�h͚5�������|�~t�Yg^~�Qx�����n�i�뮻��<����Ţy�G�iQ��8��>��J����EG}����z�U'�x�[c�[�0^xᅶK.��w/���S>t�G���_h~�c��ܹs�������2���$��r��U�VA$�ʕ+m>mg���=����}���a�4I�y�w�%�\�N8�����{  �"���ðx���Xx�]w-�߃/�˟�袋�ݒsߢ���/~����2�K�~�s睷��OAX�z�J�P:cӚ��3[M�eT��aX�:�Y�g��]�����y_Zh>��C�O���3�������y�{i�������ۿ��M��ַF�oB,�H�;�:����x͟����o^�/|�7�cKq�-B�?��>����[n���V�s�=ȶ]�
E�811�T�O�G�kS�=�����p���}��ߵ�#�M�_Yb��GWg�(֞w�9�����O[y�������%�a���i&�7����'���3�8�ܟ��'ߦ�<6;a������΃~~�y�O}����I�_���~�dSG�'�Q�t��~�_�۟�̙���t�9��KO<���7�p�?�V?�p���[�x��)8���8���E���i^s�5�~��o����1ڌc���W_�3>��;������~����W�d�!C��Ü�cvj��5Qlx�4�+Ez׻��'�x��k���eq��%�\�Cڂ�Gi�o��z���;�^���(0p�DI���QVL_��O�����f#�~`���8���{���ݱ�ڊW����5oGDF*���6zF�^W�"zz���6���S��<������k�|���?�����Rɣ�O���F+8��Htp&�f]�7,�~C�al�`�#�J柿��������AJ��S�d��XB��@N������<�0`"��R����@L����4m�1gΜ%�C�b}Bh�H��燿�c�l�6�(�_�hQ�����	��,�q�Y�����6�=���a%�f�����,�u(m��^k4�H��T��(�ʊb
����>�Z����~��G?N�q���o�Ή�MK,���Ot$Ću��j��q?&볟��������r�`y��~��w���[y ,�G����dR�_�@��,�I�:�@8I �bq����s�Y�r�i��}������?!4/��%N�f�)k(\����?8� ��9�y晃|����r�2j�h9a�t�qןq�)4oގ"B�@��⹖-?+�
i70mlݒEM	a$��d�w���ݎ>��c���_/ᏜH�a|�+_9��/���KNwB%��"�5A x�������κ�?�j�h)a<��s����{|���Z��+5�>��w�5�	b#�⍬�t�^���H@H���t��O��s��i3&�����4��$����L^��%K����vۭ5f��0.���?����B���j��ƺ%+b0Z�p��'�e2._���}�s�Y_����Q���_��'�l�$�h�����-3�[JW]}�	7�t��=�V�9E�w$���R�U)Z�`[)ל�j)a\y���$W_}��4	㩧����=�n���;f)ŴYG�)�3QA����}��ٳ��|��ߟ�{k���Yok�!o��④���Θ={6������6��ʛ�c$�����s��丆u��w���~���������`%&���"�E�'�x�Zqݖ��z�#|�p�χ��(�ٸ�b��9�ݬ�a�
�,�ŋ�e��`%o�scJ��\��w��ElOO���'''�Q�eaX��b��R܈^t�A��CصU���|;��ΫV��@<��cq�i�5[FO�����9waÆ�o!=1O7���''X�Cs�8�9s���gvn��V�X�GBo��Römѩ@�K�.ݱeץ�cƌr��`��6E�Y��&n�vp9@<��N��ݴz��Zu��^{mF��zk�D���\�r����n�k4����n���v�A	�ʳ���Y8�r�I�1���3Zu���y���	CɾM��L|D���I�ܻ����fx��&�fs�&+a ����m���B�44�u<I�8u"RxN&�����e����(��0h+�u����M���{����I<ĘDb$��y��f�ey���,:F�Di+G�y��l&�ɇ��,�Z5ZnK&hnِI�~ɢ�� ]C������G�\t8�@��c$��pQS(�b���dA��fc��|f�@�1"[[�4�AFK&�RQyE1��5���
����300H��J̈́*�O �	W�8��H�����?1<����Ds�K���2+-�}�hp����f�ϙ8��3o}c}����\=�붌0���Z�!#�-8�4���A�@8q�v�����^.��.gC���9���r��	�ɐ�$�0 =��,˥B�P�c�%�#�$
�h#��l�ha�p�+��P)�d�-�n���E��b�,�q,�cK/p�;OVrVK��q ���4�<�!�`n!��rU�pŃh'1�To�s&9��$�J����i�ò��G�iG���pY��J%l�ǜ�䵵A0�6���@�=��N�)�O���;;��B��){Z�D��g����9xUIIĕ���ʥ���N�9'��9ژt���D,�)r�J@:�E]
1�F�o ���c�Kϟo��_��;�h�5�6�`D3�T��{"�p�iӧ�?��:�5%�ϻa=�S�d��-�-�1�'@�mSM$.rȾ�����|;��|��fϞ]?��w]s���9q��xԑ�w�GN���;�8ꨣ*,\^p[�nV�8X�/��ne�F��D2�ň�Mx��t�mw�׾��2�����p���W�"	H[s`���[r Z�c���ğjU�=t�O��m7�U�t3��4>�K?vʩ���k�������~�/���}h���{�;��v?&�4+���=������7�y��@���ض#�H�8o:�pL6'W2Z�i���&k�*qpHM�G��_͋��,:v��W�.~����¯��7��v=�����8�?�o��Ƅq�㤎�5�/)�9L�n`?�tJ�D�����f�6)ul@rj�i;�/��8��aۺp�O�-�e�Ϋo�麅�v���+���/���1������ʆa�`�$u4p'�d�Ԣ�-�N�g2�|	��d���c��W	.b�h��~3�h�X��������q��_[�^��/ް�N;�:��!-�Gn�V����c`4ńZr�͇��)�dd������;�v�u?y�G?vƒ���g}�/�4o���Oc�������;bƮ�5�p�U�!�}$���%`�W�a�7w�r�/��r��xξw�}��]��/��?劯~��Oo��дz��L(��BVV�M<�8Fw+���	#����s���=������Ww���;��e��Ѭ*\��u;I8���u����%�`����1��m�}�{�\r޹�]��.�={�eW���oY������1�b���%~�@�*�?0&��1}C��'?��3>�i��?�J�6
,>v�����u�ǎ�N(����ئ�@���ͦ�~=I9��������0�/�����s�����Cl��L���PTA|�u0�ZEbu-�7%a4ڙ|�!�F�W,�0ů0�~��#�f��a��'�p��Sn���w.\x����ͯ��l֚l�)��?���%�.�a[0�:�rW�S'{M>��5y��?9s��#�Ng�V�Z��o~�۷^x�E�IE��
s��խ��shp�֪�1�6Y1��x'��~�����A����.��9p�8�1��JW�Y��c�r4��&�X�=�9F���Oj��s����s���=�<󌫘����ȡ�������<�OB���9��0��D���G�͜9s���5�;����n9s������)V3��M��F�_$DӼc3r]�b�i����}���p]�*����n{<��7�Xr�Fͮ�̥E#^7�n��[9ZKʌ%
�y�<O��bq�����M�z�u��l�o���F�VϘ��dN��m��ZB9E�1Ls�V�PEl�g��9�m��.L,@�nR�'��ko�w�̖��d�$Y��N��Y�2�2��);_�1Fw�01���Z�㴮�ũ���e˖e�I��~�'�R6��Ea�:�C��δS�7��sX�R)�OW�ߣ��[������3�<=�Ѓ�����a��0�D$�E�b�?�R�Bm��F��ߴ�%
UK��8����������k��RƧ>��k_��SN���SNy��]���o������D�*���Ȓ��0&��3�o��V��R��^uC����oe���対��Q�}�����NZ�ti��;�8nqk`j"�)s.I<�5�MǞm+[=6��e�qI�]�,tH�Q������E�_�S�Rؘ*oZ��0Y�S�_�٥���?w���y�G�������s�����b��re�` Ҕ�S��M�M�16��L.� �@nj&���d��"a跿}d��~��Z;�BVG#����Bt�i��p�����?�~�d|���G��bT�������1g�Li�500 �o�m���Z��e�]�p�%�Ă}cS��x�)���'�J��A��f�1T�WZk"������\�믿
�DU���@.{���HED5�u�*�EIh�������ъ�C�}��-�@�R���䮩�b�������A��
�a{{A��_
,&�䁠�	~?����z�>2�E�d�7e��IŜ���*��ۻV�%%�@���(��fh`܊봮p
�$/��v�$�K�'���Hg$ҟ1�j�ƍ���˚��(�0�p���5�؍��0WenL$�\���	�8��c4�1�S��jPK��~;Q�uO8�1�J���h����8���8~����`&�k�U�u�!�>�ĸ)R��c�j���)x=���uK��Vr���I1`";���̶'Al�oܦ���ٔ�k�o$z�By�ιNKJ�LF�h�WM���uG�Ҟg�>��0l�YՊ+�-���O"<�~=��U�o��#�h�Z^�>�c��Sa���cL�X�dQļ�-9�X�x���-�Veܵ� l�^����L���X��Y��Wl�h���s�d�+Y�¤s�� �N;�v2I�Os��78����
è%�d2�f����i{{�@+�;a¸������ř�>��<�(�j2Yq�o)te�\Τ�����~��ex`�6a\|��Z�j���^{�<<[���':����UW]u��>���o_�`��M��	�#�Xj;Ԩ=��pR�@d󛬣ӦN�J���B8�?����p��_�c�׹�;N`>�T$?��{<��*�-�܃|{��C���#���?���i��0C	���8�t&�/7��,�>Dzz�!�7�8�+��leSn�H�:a��$��$:���P(��Ƅ	�Z��(�b�{'�K��
�o�N o8�Ht��cpp�mS��Nr:'�� �JUBMz^�D��&`C�rH�q�R�\.	xk�4@�X��k�x���r�f�Y�(�[�2I��V��'LȎ0:�<��@:)�R�,S�M@�^_�]�1i��Ġ�F��[�ӗFI&%�L�HI��tOE��e���D�1h��1�@�J������iH�#Al ]g$����0��O�t�ϲ�U�'��1,��@L�EO�\�%����	�sM����w7����,@ {ǟ�ST�BJ���}J��3?�,N�s������HH����wS9�����\�s�ąw�YoX���&�a����&?K����D���g����#���)ND?�*�)Su��b�'�3��L�;�ǡW�S����:H���xA�`�a}B��'L�m�N�u�������2i2� ��g��d6�c��	�f�!ʘ)�{ȟ�MaP�Uf��R�n���ɷl�XS�w.��_�f�đ"�Q8F�"z,e��'�I�Q(VM����G����uV��V�R|6Bз
���xD)��a��cC��M��Z���.�X�0�`���Pd?�C��a�:���EB�O�0�8�>����l~J*��j�Sh��3x�[)?��v�ƺ��N	�gx�"^�J�L�c�x`��0�+�O\��:,�׷�I�*Lm��̘�*��e&�����:>�`̵����Z1��e��aa`x�n��i�j���<0$��P��q�S�x�@��d���ab�ۓW�2��	�e�vT�Lc�p�g�͟*g̺�W�L�$�0a\�݋�����|�s)'���Z���d���~z������_�P�^ه�"k!4�����e�[��^`���:`�[5��&ˈ�}�&Fd�S����a��hC�D�k9�m��n�F�U��2�D��,�4��BoQ�^����C_���ڔ�|���O��''c�3V�Cx�s�]{-}����ț+�`����\8���+�h=����++���������|����Ь^�����+_U�}&5^��yU�_8�4�1a�8���y|�������rՊ���N�M}���'?��<�����[�CF�Ȼ�������p/M��5cƋ/�Y]�-E:��(���ul���,5$7cF[��[4���#�X�ݫ�Z�:��k>1����V�~Xd!Ϝ!8��&Q`T*7�s*�T'����a8�N[:AնxU�-vg�R���g	1�ޠ9'��y�rW�^K�Лc��k���J�8�2���yQ*��avEp[~���o��Lyh��2�N+��]��SO>��1���ʹ"/m�N:��N��u���o���z#������&<�|⫞�5��a6���i���cPkPF�[�0l;��e�2�Y���E����~߈�]���Ӱ��(2*�遨�S,v��I��������l�a�2���A4�e�6&[6�Ҵgm�1�0n��?�;�����:u�df���%N��<6��5����AZe�������wڐ�E5��c*�����Yfª8*6�{�:n"#e�3FD���15�f��K���Ղm
�TM}������B���H%Ū�;N��xm�>V�q<�Ib��f�v=2~z��~��j�H{��^s��7�ڊ�������]uH͇�{vY��ӴE^Y<Ł�=�Rۜ ��+�� �5n�7z�7F��l�1�]z�7?������O#�/N��q[��'��s3��&��1���t�)�GFF�����(ӂɏQǣ�l����:r���L;��^s��6yٖ�ڎ���sh��������>Y��Q��m�o��T(l�m�{��]�2�,�a�ෞ�e���J`K�cID7
׍!P뇬��\ެ�N����j��/��y�5p4��>�v=��΁0GE�c�v�1-�@����۳���(�e��ݨ�{�r�Ƌ<�۴׉;0��]��H!��M{6	,����
�A�ӑ����y�в!�R�y
����:'�`k�0e�qVN�6��z8���1���9�C�
a](d�Q�Lo�V*9��08p$3Q��4����<~�i��R���*Q���M�ԫ�O�;�����l+�E��0����5>-q�����.��h�.;�`��`e�ژ[�\�VU�{��S��R�����G$�v�ܝ2�IAy��R/Q���Y�y����e�yU�8�E�De��jmE�&F.\��ڱ���pb'O|�뼉v��7�9���Z��z��[��$�a	�p���K+�Ӯs����p�������P�_O��/�ܗ�A�]Z��E��TIt6�l��l��LhU������������p㭉������yÝ�M%6��TF����ub�H��z�H5w6Kܜx8�z������,����A}�=�LEU*�j��6�9M�"�?���akǕ.�&��}l(�APhR/�G�bA��iȿR�'�=��I�=���UQ�$�A⼍A�!��x�^�F�+ejgkg��D�gH&?�K�O��(*Ih��>?�_���PY�V��o�� N]lɬ��aȵ���R��<d��L�� ������FיS֘`�8>��e
m����2��^�~�}y�u�oh�,�01��L�Q*����ג��S?�bŘC��f�cJ�0���Iq�d�m�R�F��ވ�e���(�����"�%?m���]B�(G :�	�4��g�-O�R?�%B�� �hC�7��,�l҈=F���ұ@�G�
�#0a�g�̚󹙔�����	i�0�6"��X��ux��������ƈ�2F��U=1�R��O]v̧Y�P�;�?�A�d]b5مN&��{;��NN6Es+K�PVd�V��m�_��=�}�T	ҁ\+`�� b6�z����� .'��  T?+=�g�������r)
�a&eD�j��`q�C��D���qX��+�Y`�e�XD8F�O�"-��wl�~Z�6D�2�E��&/�̈́P���N�ya��!6f:�(��Ї�7̒�`H(*�f�XBw- �d�� L�ejc%���b��/%<^�E�����KT��M7vRi96�P����ׂ�����%�ʴ��R�t
�R�qP.�F�؇�7�y&e�GT4�� JF �G�����`����+��,X4~�]���l�͗0M��K�h�&�v��)�����x��L*��>X4C�
;)�^#r�<_���o?��h`�� AVȊZ�#VH����5h"����w"�G�χK�]�Akʒ�p�y,F|�T,f�>��1���+zP�D�C�d��"�L� ���L���X;,ZB_�"�!�m���3��I��2�tA��D�
0�V�b��9EԄA25GQ8sɄ�BJG�� ��e�?�)�J�]�����X"�J��|QF-��.�j���0D$�S>/�
>�7d!Գ(U�l,�0�J�r@��<bšDgRt3�����q�r�M�F�T����[�S��V��;�&%n���6���Ĉ���G��^4yc�Ԉ��6�$���(�6-�\H'�p��P�
�MWēMUb ����WFT$��m=m6>D_/䟞(%���D�Hq9C�|%>#э�rMj��P�91�y���#���{C�Ew
c��"�_���ޘ��|���3R8E�(�.�Cs:\_�|Yej��cXcG
3�5�Dk��^djq����;�R%��0�ݑ(�"!��9��P���'�D�C��W�/�J_��{$�(9���,�G$,�l&�	W?T�b�sX��
y�9e�B�
�iQB��}�ܲ��`��1��Q}O��8�|���(�0�c�F��(W��:5�Zdَbq��WT�v�T}�g��}@/*`G�՛Ĳ4ʊ��Uiu�;p��5C�e��D�	X�����	&��(9��f��p�^�H+�X�HqAc��J��4��v��H�[�8�1��>�d�����G�m�,�S�u'�>b�����BP�q}�R�5SDф�|V���x�.j�#6�M-�#q�Í��F��5�U�]�+�M�/L&(1g�������������X�bs.L)	����(�b7�[�2��B�ն�;��w�S$�Ѱ��~�h�T�,��<�Ta�_�
�{SX����8 n~����7#�,d(�4�h�4ŬS;
[�����xN3���"�E��j�ǉ�9�a��8Ƹn�(pvf��7�T�b���Q�Y�ld)U�PրUi�Y���bd�1��8���x��q�k(=A�%W�.N�9@鸇��6��6�H�~"1_�=\���&�и6a@y��3�\l��&��GyT%42��`�q0ڢ!�`]�b�ITi��xp�0O%�n��[X��Ӵ�G8m�1��q��NciKqb����	c\#VR���@�66��g�����O�� ea�D�(d��q�dL�K�&����/>���b�6s��J�T��UWe #��w�*�v�4d�4e%4N�F��L	���XU뺎��*:1�� g���i�h�9Hy��sfQ��$`�cS��aJ<@�a�邖���%bK�h�ڃ5��5��X�-�s�����#�g�Y�0aq7�{&0 I6N�8�bļ�,Y �f�E�B৞�z�Q��t�OJ�Mg�Ao`����Y��<�ê� ���������Ar��^��!�� ��'mJ����2q���sT�2�@��K����(�-��9�	,,�D��4k�:�<�2�4��I��< �: 8sr���T3�;�c����fnQ���i�[}�e����"B�j���w�b��mJ,V=;�&{�Z�Mִ�@F8�R=�aċ��J�.S�]y~�6f�i������W'7��)S�O��DQ���m�PDQ���xd;���xK��d��A?�d�����+N$J_�(Fù���P��fã;�!q!'��������H�O�Kވ��"T=�JL����
|_&p+�'+,�����aQY��?��3���+�e��,X���O4�ﻶ8�&:�h�$��W�'ɤ���9�M�ޫ�rh�e�c�H��H$�XIq�b#��0qYQo LS+ ߫0����+�H�Xs'^�����e�\Wi9��i���I�E���$M��	8�T�8���F��� �jHWg��Qۜ�C���"��:�ق�Ļ�(mz���ɅŐ%J9��L��e+/0�ϊ<b����	�X(s�1R�g���$FICX1���@�c��,�W���=}T(��*�F�
��,o��� �j�)�0��1�ɫiժ�|BJb� �������R���7�o��Z{� �IT���$�u!6I���Sy�^[��A4��K��1qx�:�9C/K��	ϟbQ�fh�LY�2_�.��:�N���(�#�f�N3����>�Hq�!Kt�(gieSG*C�ę���@,�b�����,�"�&�cK��F����UQe��㇅�Jj-���;�#�Y����W(�1A�9*ȸ)����;h(J�uR��X_�q����wS;�D�h$!oڀs*`�XW�5����l����O��sur&���Rm4�{��,�||��2hwQ��x>X�j��!�'�A��J�T*�y&�
�_�bT�c6�� J��1�'Fb�Xm�#*� /@�����4C^,�x9,V:�[%yRBA��X����	��Z�,k�a�5r�a����]1a���ڌ�tl'A<���iPܘ��}��t"Oղi0.(���q���!$y�E&�
s7q剗��P�]��\�N�_�����N��>d��C�X�*���� �o��&�Ԭ=���YN�<v�I"ǋ�:ZL.�j7j��m1�P��7S�6�S���r9��g&d���Krt�z�-`B>M��i����/1q�
��f��9֮s�Q�aa��FcP�L�����s<ǩ"&�&]�V�C�R3i��Aui�w��$��_�TYl�G�%L��c�e�N�)����}�,> �)��0��z!RO��56QbF�V@��i�1'OE֜ײ������s���ryuX��]_��ꄋ���^���*�;�l۲��>E=QAN[��XD �v����(�ǒ9��9��N	H�CQJ��<���F���	Ew	"�1aDl��R���Y�xc#�Zz�.�]L�Y����{2W�dR��fѐ�c������k�#�ֳh�W��Úc��G��D�&쨋��h=ǈt��j��)��Yc��'ކYa��~����L�U���@S��.3G���8iz%��o�	Wx+QM�O�9��Ma�s! }"�P���	#�,[��\
�T��"�Ֆ���32$Fo����x7S:��f"B#��b���u��>�F�:EA�0 ��u� )����(����U�_N�oX�QJ+��j=d��#��ۈ*�ߘ��U51��ŏ���2J�K�������ʬj��M�I�\�I���F .���zVEW��H]�H�F1��]��j�Ni��u�GM!�
b�/	T�U棸J,
ewF�x/Ԡg�pr�MQ�~���§��8u�W>�H=h(1I�B2��b�a�U�C!���0�8��L��= L=��5��&J�5��G	�N���t�ر������2���c
�K��]�K%)����^���rRH.S�bI��aE�"��Dj�L|�����Ig�ћ$M"V�6��� 55Ľ�Xob<B���3�1�B�u��g�5R�	_j��G#3���&!*xK��c�J4�h����$�@�{_��u���RJD�<�OLlDԌAR�K�B��j#"Smr�)4~.�HGx�i�@L�d�k�i����e����hXE�Òg�@#��"3�֐�`���¶N۰5��z�T>73�HF�s$�������J94����������a�a�cWU�� CgV�-�G�hK����6�c��9'��ǖ�M𼂫h�7�Ok�(C�.�M�Ex�r�)`��TF�4D!A���Ñ2UVL���%�BHEmC�)�J$vMPǰ���ݫج��vA`�á"- Ԃ�fɡV��u�-Pe>�B�x�n.�xf��@e�+(P�;��fJ`"B*��RJ���R�l�&z���@����:J�]�~}E4��E�w��|&U�-��s�Ɏ96D۬�$6��]�la�n��%2U��V��g�d��H��,Ca.BC��f�'p���@R��Vk5�]^ac�K�/�7��4C��" �%b�R1QD.��&���r=��|�8#�l��gR>[sE�Fl���:�9��G�ceu�C�� b-zH�*F���'��6	�3��6��uٮ���H>����QO����OB�tq�H@>��T|�]b�=��Q�[��K	�R���~C�Vt�0)3I�Y���ua+.c4�9��G��H/�Dt$�*��<�5	?�!bn���5��'�X�0�cC�������_]��U]JB��Pu*��'�~�ծ�C���C%*2���i�s�CQ�Ė��W of
KV-Q\-����g��p��@��P5�ee��بD#h`*c��K��Td�P"I<��b��\���馩ce(���U��YA��6�Y�9Y������r�� ��^�\�@�rI�c]Х�����t���|��m�i�	�75�GV<"�m��)R#3�K�xQw�;�-��������L�Hsg̢:9�3R�R�����ry�"��T;��p'^NW)���i�c�!{���w��uk������U��Ux�r�i�P7��c�)��ԙs9)�x��ixs��>�r�5��|�,���bţ0�Pn.[ ��VA
e�Y�dޥ��\�t�]\�N&+DЖM���NTJdY���Di�ζv���g�à��6�_ˇ���*���`�*�%�I�����ja�	cc�.I�x�b�Lg|?z�e�'�7P
������Y9{�fP��3�|ǟ��/�P��)���R�r�H��}팝��K3�6+ǚŮ���]������3�U�pTS�\*נx����R.��b�`�S:;��,xa8|��^@պ'Չ�s�Z�*��(�L�" �2b�gsm�;��5R���4���V���LA���v*R.D晋Ʈ4P*Q���JuO�7��2�<g�#�B*b��զ&��h=�����% `�o�#́�/jh.��57<G�y�L~o��3��3OڃY:@�W=A5�sYތH�Oc�&��A����e�Sɢ�5͞Ӭ��i��i4��#�u��D��5��L�u��a�`������6�������I�:�;�8T��y��������=��C]S
⓱b��������S-ɯ�T��ďA�j�ژ�Qq-�S̩�}�N>VS��w����+��)�E�P�Z�klvQҌ��U���T(�,>P�J�b�O@%v�hM�F��<
m�=����]��󎦽:��������Oh�L�����f*�]s�3��&N���g�C���V3[�@�4�4E�_�5����7���1�{��Ī�ۦS�u�����wҒ����;�F�z����^�ǖ,�߬�:+�(�]G@�Jo{�|�6�[�R���2�˫=��s���A����6��޵�n4�};Z��rzt�2ZSdn6c��F:�s�Ϗ>H��:�FE#Cw?��E^A��b�*9�/eM���;�=�@��	c>�2��$�2LV���cy�tC˱� wb�O5!Y�ev�V��%ϧ.6W�t,q���{�dyfO�z����TH���נR��U����B�$z�L��^��v���o{����_,"�0��2��3��ϡ}�a�Δ��Υ��w.�{�誟�KSXtt�N�s�NL5W�m>辍n[���0K�t�>�h�;�q��4�Ŝ飴]t�r���%T��m;��>w�,�ޟK'��?���h{�]�ɺ��}�mM�DԢ��K��C�jLS�X�o��u1�sR��xuCխ�ݩ��P����Þ����O=K�f�@eF
��TDَ<�q�+��_�N�6�˶���n�1+��n�~��(CCk_�?s<��D��@O/]EUՍ?L;���^T��*Ma֎�co�=EG��m������S[@�ٓ���K�����N#�+g|���O'��jƌ<�Ȁf���`G�&�Ǘ�x��.Ru���}���鵥���DN�j��D�ͫ�D�|��5�)�1���'&�%��8Nb��T�e6��gd�c�Cec'�J��.E�L�WV��j��rJU�>�߼�������މ���V��T���Ot�^�U+ג��A��p31�����=����)8��t��t����>���|���_)�wSG[��Ţg]A/��Y*t�(Up������Bއ����Rɤ���G��ȓ�ߖ�~�`���=w������~�`0my�ӦvRƝFC3�r]�T+�N:R�q��p;���g�a���.��t��С{̡�|��W6�7����>�gr;w��U@�6[=�H$Ш�P�D_Z^e���h����H<��M���T���c&c�-rT_��,>}#���K'���t���oK����CV�2)��E�jm�X"��&�,��;�?��~������_!�}Gr]��̻aV�	�urbjZ�n��g��wn5h�C���}|;�cv�~��g�}j�fg���:���O� /��"Ųf��X`���=g������&������W���<��{������˾y
=�2s�_<NO=��ܮn��Y9�E��{eo?��S%9{���K˗	G�u�)R��ηK��g_x���v&��L�
�$�}�e�R�*	��;Q�vC�j�nc�4GUhA����C<�JG�y�$�ꬿ1�Jƍ���Nk�B��O��=_��6Ņ�*��zY�ɰY����>�	H������}����NL�_�yz�Q�Ko���A��LA�TI�R��葕颊��H�m����u}�����L�;�$č�zm�z�dQ�Γ_���ZCKW������f�B\b��������VV�}�ܛh���л�K��>��g���C=���)}}��Nz�C�C},��R��M�*���YJg34X,��`�:��"+�[gp�	�(�E�P�W�!�C�FO��=�Di�����,�H�(���[_i�[@���]�3R���VO�
�%��03���̲1i�tɝ:�V+���W�>���nt����1�?�[j�兒�5Xe��k�f��YNէ뮿��z�I4�Z��2)F��*��7�G~��t�G����ffS-T�.L�[W&�Jp���8)�'�*�*�f3a9y���ӭ�Wҭ����oٖ.:k�y��韮�9��uLgQӖ�� �M݆*}EVZۉi� @�V�؄-I�:9<�+�XgE<�fn���W��Т[��ſj8B$k�u�*cH삂��m)���@"k,e������g!,��_<a*�'��)��&"nqKN��e%U1���z�CA�ewz:���􁃷�SNؙ~��+R�=9�٬@�C��U�y����֮RT��>�@��˯��5��5D{�-��c��S{�@��O�7{6E�L9�(Y)��&��,[E�j/�Cm�5[(��@Zߚ54���?��O=F=����N�V3Kx�W��mK��so�颧�(W���#=PD�ݿ{�RLxq�� /W���1��L$�C>����pB1�"��L����R�0��4
.j�b��0b�{A���oF�['�W"8�並�*�@$�t2L �����L�G�Iz�C��R���H����|�?[����˶��7<E�|��t�GХW�GS�fP=����Ot�ns�c����DԻf�,����=w1��'�0�X�L�MW��t������s��ޗ�^�mfmO;��AW^�$�i�R>}3�d�Q-����T��9�O���Y;����h�w��I䱂�ڒ?S�����hG�W��˄m�ѿ�F��mK��z˜����>Ms�sz�M�����WXL�ie����X� bf��0'AV�ҋ�fPcˌ���d$Y=*4���*a�t<%��a��.�k)�16s5�6ݏ�S����$)EGU��zN�i� ѫ��t2�~z
=����f��LTO�iy碷�n��l.�؆�eJ�w�@�����
�|�4�f�c[*��'���_��=�2��N�ryz�%t��K���^:�sD4�ġ��Ѳ���A��
���Y})��ζ.�f���f���c��N9r�cޮ��S�_K�_��D����,�"Χ�^r}����C����'�f�r��k��w>Jv���c�;OO� Zœ�����S�4"�ď�RcV����ƪ4�I&���^(d�ш�*���!�	����F�%E	�3�S����.��`
T�M��s�J6���`��ѓ���w/b{{;�U�6���x�T������28eZ7[Lrn���֣~���L������`����g��B��V�C�C����=�)���W�be�����P��K��U�εI���`���^���>��{�k�j�nz`�tσ��D��NQ�Q��]X5�K��k��ϟ��n7���*��<�X2 �e����^��K^�+���ɢ�g_�;R ��JRyQx�(��.����+�N2O�hbH��e������p�&����g�~A�L���� �����S�PQWVP���uH�j�/	�>@	Hf��w���Q�!h�Fqp�P��FTc�5t;�$!��i�WA
CPS����)TD�8+���`_ޜ���b�L��,6��J	'B�ӻ����_���i;�[G���HY�q2�C�mn�#P��$�XJO�#��k,G>����p�Ä���!��ܬ�d �{K��b�l��3V����4x(�b�O���aB��Gg�t����@��q�p��o�v/�k"�
�S���ME9�5/}_`.���B��À	�C�'9]"�,S����P�[ .*�,-m
���*�WbK()m���A�=�m�+b�s��B`{��Ҩ�㤔R͛�+�F�g?	3�����������
Ѻ��<�X�%��B(=���ʉba�l�j�l]��a����*.p�=c���Y�'&VR�-䚘�n�
,���_�V�RA�H}2�GUAccI Nc!��U��G�e��J@��7�AJ?M�O�@���T=T�A��T
EN|i!)�Qc��P7(.����Cĕ)�{2�Ȗ������n��Mq/��#�%a��s1���"���b��(�^�RU��������� ��!PB�-��,Sk�MJ��!�rb�5' ��p�T�J����Zj����G�A[���yҗ�?���QT�ut5�WY|�'�<��/�k;��0�y1@��U�S���wL��NDo9a[�п��yA�@��*a9�eE�/R��Q����X�6�t"g�)Ś���V��/�`��'R�l$ʲI�Y^ &D�!@8 Ѡ{uʲ�$ռX
Jy���l��5\�y���8�R@N��8�9(Ub��3�V����0��t�s�
��d�mR����8�XԘn�P��V��51E�Y�x�� ��͵���<�����T
]Ή��pe]��]pٔ�P�֕ �X<�K���<���(
�b���yUI�����C� 5��U���	`�+tba��	��v�R�+��,��eQ���	��h��I��@�����ErA�<�j��rA<ӑT��-&$p+�l�.��M: �D.��1� ���LmF�C���!��݉�`���	��@8�ͬޯ�s�r��t@2T��@O��a�5 �
O�*�T����e3қb�R~X1��@2oul��\>��t#I�,y�A��٬bV�PJ���׵�(��6{FG�8Y9ˣ�W�P��*�_���f҂R
�jC�h� ����8�N�ιT���IʋfI�;X�S`�Pz�E�{��L&(xUQ|%��*W� !@�\p� �w6!�)����s1,0�[&B�yl+�,����Tx��[$Y�!0���y}͛
L)����!g�n������,:@U�O�*}+�//�bsHǄ��e̛��k�G���*��<Wg:M�>�� R����gB˸!�X'q��4��%�mTS�@w|B�^�s]�H}Op|��v�ڶ��(�Tc=��=��1J��1���U#��+7^I�Dk���$`(]@C��A$�
�w4��mw��Ա��T\�Q�*$������釩��Ս�0�+T�.��U�V�-�l!̢]�؎��4Q! .^�s��O�-�5��x?��TH�*u�G���z�#s�&;�N����̳V�����]�C/>��'���ST�~K圲|ϰ�8F5u}��#p�}h��?C%t(w��D�c"��x���??I�������v�K���!uN��5P��/���?w!��n�i�������A�o���@���g~��e�����(�0XT��-�4��L&G�����IauP���l�y�!�A�'�v�9��y���
��{���B��N�QřT�'�レW������_,�c����\CJ&�L�Pl��#^�iوf�;�v�1�Y�R��k��9�)���Eǭ��AO,롔W!�S��<s�|�u���\L��wo:e���5m�A�ʞ�,��3Xl�T�n��b���s��l���e��0���Ru�������fNTa�H�/b��h�DA.27~�5t�od�X�����'}�bS�3"~�'��1�5�E��\���6D�n,09'@[&պ
� �D4��giv;��� �Ѽ�	�w�芹�O!��Q[.m�������󑥓yP#�9�\�)Lp]i���*���7|D)E�;�i�	������+�E��iR��Y�E
���H~2���x���# i*�ZET{����M{��Ւ������b���b��כ��� n���q!��q�c�YA.�/�k���^#�Q#ҡt�cBj��F���*K��|�����pC�Ft���kؔ�H꧅��}��iC�e�uO��@�fٌ�E�2��{6��rq���4���3a��|���AJB�p �ԅ�&f�_3���&I���9�p�C�ur"#V�Z�� rB���$B�H�M�	���TX������%׍'u�F=P�bCu0lG5�&�R�R�M�+����q��|�8Pu� f��bԓ����F!:D��y�9N�)����
U44�k���5���yD��bh��-�_��÷�z��Q���~ �lE�ե�)C&�H7��m 6���cH G��(�v��L���-~~P$��R�����n�@��sǺ�f$VNzv�=���4t���2Y�W ��#
!kZ�����bV��L�)1W�r�4BK����gJ��##����瘽{��=� _��-���T�3y$���`H?�x�j]�d�\Z���J<��T�*�L�_I���t.��1p�2��=ߴ.�y����etKJ���{�:�M�Yʁ��߈Ԏ	<ޤf&�� l�*���}�ڵ�7����F��]�d@6By��,�8#�k8�$0��,�\I�'�(p�pU�$����K�Z�|���Hm8E)J�d�Rg�@�#I@B<:���T�"!vd���ä��@�Ռ���
C����J ��b*M�:��T�@E��GWrz-d��򘉠�x�̭`���)I 5?���Q�IٮqA��[8�Ⰱw�y'-^t�,8F6�j�~��E����˧�$�9m]$o��p�.^�.���
���:f ��iB�C�It���ZU�P`�H�_��T𹧞x�.|�/��N�J��}dQxA+v�WgQ�1�\ fE� .��"�^��sK�H�ܼ��H&rTsa$U�	�b
��z��]Ya1���Ɛ1\�UED#���(�?��ZJ�C��tEUX>lt�d��M��\P³&Y�9o�����5��%�!<�._Nk�RcS���q�r͆	
�){���]��c7Q�g��Q����^~��[Ջ��\%��~�4.��F,7|��R!2��¢�� �4ܲe�؊,�e��9� �NA�����i�+�C�T�PA�j|(�lGC�����ء����]R0=f��w��(��দ����a��Ǥ�[�,��T�$�Wzı���֧�s(�h�ƕ{`�c�ch}e�S���/7���C÷�:�&i!jd#`%�I}��l"�憱�!l|����7��-uC��b�I)�O)g���M��i�?��u95�>r�x��-�v7gش���t�q�aȦ&!p)0N� 7 ��=G7߷f8�~�ah�/8�'�8���~U��P}\��bC��J`Ѫ�}t��h]
i��n�f6,�&|�F�HQ2�lwY�jU60�\uBI���.RM[�H��}�D̤R���e��ͷO^�̵f�1��IZ����{:�3Ho�с>(���@�MD�noXA��'=�M�8<GC+¢�e�&�,4�Q��U,�()����d�|H��@�tD�F&Y�h���EJƽ./)nR)P��zS:Gi���T���b���+�F�
$��G%"{�j5N�p�X�G�ԼF^/f�����hː,r�g$'�AZ�l���=4T_5�u'�l���9�b%�ћ,�cP��O��zC)��q��M�Xx-�H��b��*�I\+�8,5��~*��V�VR�]B�Y�YI4�~����'8ҏ�DY�.����DJ���N=���L��Xz$l]m*563�UJ���aqE��d��6�q�Z��78�*����5�&�����Ł�:�(D��'�o�������:����A(�X��$��֩���br;�5G��i�u�HS�DFb�V�+)�I!�ULE\|r�tbQ�j�XR�Η�R��A���]R����|n�\�kl�jQ� wx�MK��_���F�"��Hİ�qZ�L]K'V�U~���|�:���0��Oƨ�����olA��S�E�tm��X�%f2D�IM�XNw�X���0�D�$AB�����7)
&iAb͑٤�5�X�r�H�q�J�׎�EL#=.ɻj��O<��-BE�5�'�
bڊ�%��F����b��0�M��#H8���/z2�eS�8N乮5ּß3�T��M;���Z8ĉ&@�@b�(����Nn�7^b=ڿ�|�GҬ���$��\�x	Qp������Es&���Yqn�|�5"�r�?#J��@�,�z[��@�Z
*a(΀^1D|F{mEq�_ƺy!� Z�|����4�Q��x��{��ـ��3}M�\�ډ���xƖԝ�8@�eDB�]�E��<)&�>�&�$Wץt:K�(%#���$nr��f?�'M����:�ǆ�a�s���~�+�r��ZO&�����M����D4��������f�~mD�%lisyx>�k8I�ў�X1��F��9#)�/(�f#"�ՒI��A��-5��X��5���ؔ��:I��Γ�=*b8!۳��L����bSߔX�/��0󖕇|�~뇆����8(3W~*�qC�S������3����[h��o�nh�=)��?D_}�K�S��Bۡ2���+V�A�5���[��W.ن����UOc �3���W �4��j������ت�$��_mW���'($g�hY��y�9��o"t����R,�u5m���l��wI��ύ�(��I�l)t�����I�H��:�ee�����q��rP$y5���>��8C!�%�,�7ְ�8P��Ke�cO���/^F�G�Uy���"�,�f�T���}������]��Im!I�������G�%UC�Ԙ �� �y1~��o�k��{2kub&�����Z�i��ZV��q.}���yC��	tP�L��� ذ�.ʼ���~�a����ӨR.�:&�~U�8W��+#e��������c`�D�2�Q�X���^we���G��:���t>h6^"�����3im� �ӷ/��D~����R;Rj�1a�wHFv��M��CC�(P��q��d��j&�Y*JP-A��A2U�����Te"�{��l�[ �:R�q�LS��-rR����s(䲴��QP#_��
^�z/�S
4��ç^�fT�&C�
b�/�@��K锋lR�yS�  �Ђ
���󔚳-}���h�\�t�cD�+�ӓ0�}O�@��8ڼq�.�o(�d�am����>�)ʙ��³	�#P�}�Ȧ]�Y�:����ԙ�P S@�i��zdk����#���qX%�+�@R����X��)}D�TֽPp��ՙ}cC0$�� �a�^�veG*�!kCu���Q�>M���-1� bº�<٬
�#��Uw�$�\E 4\�m�.p����!�P�sF2S�l��<�"��Yǔ؋�Ĉ���r֘;����$5Da�tB%j��d��=�|���I-H��*�-�n�z[D�� �Y���C�ֆE&�Z�����5�Ni��@�!pB�ZC74�z'	ϛ�*��V�T\��>�S
3�UA���
��)���Y� �am:���E6�Do�q�8l ,�i�]��a��, �ZI-	K�X��Ѵ]�y��{�U?�5�c�*/�a��Î��c	9�ir�4���(#�<�J�R���YY&B�9+�U�k�G��7�j(�r�(џ�������6�"T��+��"E��G�H����%�2HE$�7�xk���6`"o�0�[#ͺ9���2y)��0t��ʴ�Z�x����](�	������e)�e�Hl�Ʈ '��,VA
��Ϙɦ��pr �N��&�j| IP|� �C����AҸ�HR�IԵ�@��㴊^�VH��H� 3pS�/�X��r��{rr$����h�R~/a��H����\L[~5T:�'�A�JAL�ؒ�&X]Et�W���`��A;ɿ1�x� �Κi`�jŊ���{�[�U��
;�*Wu��PMGRC+ �(�p�>�
"���lT�\L�- ���%�D��n�s���\'���s��ϩSU�T5��}��+v�s�^{�9�s��? 6P���{������j4e
�� Gd��zm��tݼn�t���[@�.i)q6�0R��ܥ���	�Mم#m"�@�:+^C�xl����2!�����ma̜����J�,`,GS"��5� �\l����u��! W�\B�0�e�}"�p$���1HR�E�a�vN������H��S�o�R�A�K���d��bcЛ!��������إ�d����5,e=٫m��z\�ְ^_%��5�l-\���We�#|����O��2añz�\�
�S��p���VD��J�b;���v�u1�F5�,���J>�wi�BS�f�X��!���u�^(�U��He!�q�\�\����b�¡�߹J�m�AD����H�n4����v�Fq]��~o���6F��P�����������gMT~��螰{=�v>H{i�����{䋍��)<��/�6�d.�OCTkl�0�����g��U��}��U�Zް׌l`e����'�"��ᨅ�v�x�-\�l����#+�	����Ae���ρ�!�(Ҧ�����p���H桫;�R�nӊv��d�<�����L���+���%�XT����%?��=J�=+�<�K���I�F'�k/+�v�U��9��6?��}�Zg�*��[Q`�La�XeA;`O/V���U�;*yttȩ�q�/]!��U�"���tG��/Z ��@&BW�3��|9���Q�B_�F�-��X�Ќid�������2,O�.�!w�K�A�X]bd�Kaf#�ʀR��!�B*цQ6��q��ܴ0 t��U�A�:A�� �fcQX4�����)pH6Q���Y���y�]��i��.Ϣ��f* �nL-�v�%�]��ZMVJ����T�����l�,.LmC�,�'wQI��FS��_�8c��^Vny�Y�RL�GDAe�i5�5�W����p�0ϲ�<)̂���`��et��� 4J�><�1,	�6��)Ѐ��+>0s,���B�Y�m:AQuq��w��yV�oҎ�»i��*�`�vE0��'�ob�@����+-����"��L����H:F�_�"��mjC��\�{[�	��s=j�LG�!�BZx�z��8IՅ����.���Պ�]T��Ŭ9�ՙ��υ�}&����j��)�s��	(��UXw ��yMթ���؁μ�,i��PP���16���Za��U���X��������+���M]����(�o�pK�z_8�Z(åp�8<2��ƁұN4'{�_��)��ܒ��z��͒.�B��#S-I}��al��|�ν�

�͊��/8_�H[��.��>�,qU,��k7�3�Z��k�l�؄2�`H[�B��,k��y��T5AE@_'���I��m����	5zi��Н�Y1��3#
���<��f�F�}�;��L�����8�ź
8��C�ݑ��pz�b'���Zp���3o���[���1*����<F����-\f�}/�@εF%�Mb#� uc��}X��ݷ
�.D`5!�������G�\~�:��8�q���P�h�k5�.t�[>4��Ѣ��otR�s�	P��깎� {1���s_�,1NRY�s�ե�8���u� 3��֪����.SF���zt=�%*"v��PP�{�Ư(��5qWݼs$a�,集
,�P!��K�ّlKo����4��Y�gӧ�Wg���K����T>�3~|R~�ޫ��0�Q��XN ��˂�Gi�-97ͱ[h�U���`ߏ�j�	DY]f0>�&�XPL���\�AI�� ��|�C�|�v�Y .T�{�����[��Z�w���pж������5p��l��✹��Zs�9,r��!g|�
��7v�T�q�[H<�׀%�Giuu��PL(�TG�vY1�tn�,׶ �5w6�-1��q��~���7�n�=A���]�ɰ�%�UQL��?��ی[��������D���wcY��E7e�n�Ge��TaƲ�쮪t����:C6��J5hf�N5��@�����ӻ��j#4�5LF�wzd�w��r�Li�̭���`"�{鉱��(\ř~6T?�` ���**�V?��ĥ:�X%k q:kU�;}ͼ�Z������HS����}ZGr��!Υh�u�l�$YҬ%� �l��F�DE"���
��L.��X���@�x`�af���<�>�h����`�ff?�����A6t�^U�$
,:�e���a&x9L���bh�
��/�Ԡ��c�2���:�Y�`A�9��/��$a��硆l#n�2*�r��瞑ZX Q��QW�Y>�<�`�A�nQ�UH=Gܥ#��Q3bx�:��I���*�D��պL�����D���P�N�-��6�j�g����b\.��ws��2]�x�C�p�D�����C�G��%��pp�v^�8�yO�7��
0�la�]���!��Z��0C�x�WG�P���D�I��>��a%0��Tpa6���j:�қ���<�s/C�3��x���J�|�g�>s�΁!�C��~���}"��� u�-�)f0��`��X�1V3EH^W���Şu���ݕa��IbB��w�^�EB8��P�6ѐ��;�W�D�z��$�A72�@4Ks�z�|my�����Jn���%�����!�4!���WZ8(��iny�^�D�ZD���Yw���u����JS�� !�U"cĬ+mm�.��R	�
J
gZd��-3r
e4�4
�g�<!q���,���0�%.��dlTDd4���P����������P3�)Q�������j��������/w�F��6��?��r���b�G�%��l����`K$�I��eW�����\��7������������!�|;�>�v_���|�&.���!AA̼�l�O���%z$ϥ;L�Zv��t�V	���KQg�,�(��T
�\̾�y���~#�'�Z.[��W}6m�6�sM˻ ]
;+�@��
�}��f�9�f�G�j��1&�A���
4>�:�>�tSm�^q�B7+u��^p�mw�o��>Te�eH_5u�,^���zo�B(�bb���;����mh$�)4-�܋g�}�F�T�$*.��ۡN�W��-���,��.��Y�*v�y�\��
9��ݻ8ğ���0-����i#̓d6d�YS��Q�Q��w�43T��<-�{V�x���"DY�����OGd�q�0`�42���������Q4����ް��~������ŉU�m� ��pWDJ�ߎ٪��\U� 5:&�����T�a&i�Ҙ
/��̶���z�E�����~b4��/�E�Wg�R)_�ٛ+���5�C�7�ό�شc
�c&C�����Ǚ�6�s�U�E���2�-���aT��k(GU����'��T��F�`�o|��ȿ�Ux$3\�9&J劓����>�pn�]�	ga�1D ���9��N,��	>�8��HW��*�}�,�|�`��W�m�O�Xl��3 �bע��}�f�r���+�0�@��͊,L����{r�K2�K ��c���i1";�i����-/C�N�ZB���-9�d]Qrj�2�9N�&�H��̊���=�ϵ�4W��X+�G���0%�ݨO�{�n�v��6��#�in��$��5(
�?r���쇻H���E���1T>���Ԙ,�����6�g]!��}t������|O���Υ,�!��xJ-@5�"�*ɮ�z�+���'�S0ږ�΁½$��՛.f�3���"{C��I�B�}�>�X��ϋ��`h�ܣ��E�
�/h0�р��QXÒ,��K_�2[�>h�7�Uq�D[���l4�:�Z���ܠ�!F(�B����=����7��n��;�F����zzSvZ����fw���M���0L�T���Ȫ�#K���j�3��f��v��ڝ��wYp�G

6��c	� ��7d����^WR��2�hN͡GHC�����E0,��ʼ�US��(������5F�סU��R�)�
�X���*e�(_N�b�0f4.�>���Tm�HIIe���Нi^��M��&[���ɟך��~�\��w�Ei-��i��k���Sb�,n�<���F�sT���w��-�$�f1��s��4 �tM�Rr��b$uW����*��|��iw-���.�Ϋ�
��&��:53'�`�p2u�%#�!������ה��P���ke`�Kj�2��n����a�C��,�%�J
p�!u�W��P�$tY[U �Hw>^�cÓ������0�B�M�o�>	.�1��ݾO��!`� �1L�P�0\ڨ��r��ah�AUl"�ϒj�v�u1ִ��`=G/Z��f�����0�0��K�Q#�Q�ѓ�C��@��}:�=b��	�Y��\f+�Wt:��0�PC4좑�P4�p�Tu����,��@p͚�ϑ���a��r�n�|j�Vj^�>�X]0��T�;	]��ik����;�:�p9�xB�qu��C�'�Da�պ�0FCw�裨�������	��x%6B��ev Z�뿎Żn�x	��>tn��y��X諺U�0��ynGq����ð�I1��;o�[���Z��j�Lե�s,�9}|�C�ð�F��*�{�s�Q�j���7X������׿���[s<[<�w�󝘒3T�?�Y6�Q��� W���݊~�t��#?����)���(\8��' �b�Z���s�v�DMͤ>��3�)�q�h�5�F]��p�5�B[dՄ�zwӒ�#c�ӊqt_KTv�O��v��ۀ� 6��\O����-c<�5aF�GVm
�[�c4b�E_��W��K�ߊ>P�G��=���W�0�5��nY���Pc�I�d�k�{�]s�w5��[���'?����"��������ǩ��0+��6Q�fk���5�a�qQ��%�&8��c!�o��@	N�1I'!/W��(lyc�Q�<K���^'=68H�qA�B~���0���ep�
d�Պ%ȝ!�X>��i	�Iu	��2����G����MEgD�g�A%�L���#�b('�,?�C�x\oԔ[�%o�LfM/��g�NL$�W� o����F�F-W��A����z�P�����:�CW8��'�l��ԁ��p[��ŧ��1��,7�f>W���J��J0a��i�c0_��p�9\3h`1w2��/��X��Ɛ��!�e������G�����͉�E���\�z<��;��� Y�2L����<`3��+��+]ݴ��n�s1~Vj&���BSs�D:���� ��!��"��D{Ք���+y�ۑ�H��X�4PF��A^X'��OF�$�(���9��rNj�ɲF��^���a�,L��>sJ�\%>�6���H�Pj+~�J��-\J8��s�*�d*����!{lt���$T��d,�K�����v&�n��R�Z."�Mt?X����\^&���5bEV��H��G�T/#�ˣ�O��c<��h�m�-��lsЩ,�
|
��N}��qҞ�\V��F-�v������F�%,C)�j+���tz_�s����E��=��R�j�0S�si��l�[4��eyc?���Zv�%y����l�0i�\�Y%����p�ى��^��uW&���3����m4�Se4d��j��r��\�ء����׮���������XHá��W��9��r�3b�u�7~@ꈀ��U�s�p����i��3�z-���\�F%����Hܢ�(�W�ԹID���$0ʊ�0�Ct�*6?c6�V?jq�����䮖�ԁ��y�P{�QrG儮f5O�jy�8?����劣�cC|ٟ�/��V��u��:�YK�4���p�d������B��b�����zf���>��3�׺������h�lҠ^��f�S���*Vh��C]dj���!,,�Ccj��h�kDXL�$�z��=�Z�J[	w�K��P���]��13�p�uX8�X,���+wlP��`�Z���X�xbT�:b���a�bLD �a��'�@ֶ�z��6Xոb|wĀ'�wsfN�K�b����Q�k?�#�[��[��.�$��F�k���Z��`�#�� �O��fU�b�V����O��d��M8���H��X٢���f�J�#N��B�ZeZ���μ�"T�ieVL���Q�0��=�����D��AY%cS��A��P�S�qR��5�ﰿ�ܪ�iH�=�B��3��W��/*�͋�ُ{���oV��[�0�q'6nݩU�D�ٲu;��E�sF�Q��Ë��Cp��3l�n����a�����X�N��R��q�]D�]¶3��h�u5<��޽���_�+x���e�y�h9^f[b��p�w���}����s�05C(��QmlG_��bs�Y��Z35�����>Pv"c�����������`����'5�5k���{�`��p�����?���6�U�%.�d��G�.QwX��*��X,����{�w����;о�غ�Q�u�` ڦ֘B��]|�Y$b�(~W	}ߌS�$�50��*K�h��٬e��Cr�����2�ۮ�]����ڌj��ޔ܁ͧ��FA��p�9���5�Hs��o��G����5��3�}݀Ab-�A�2����$���G�	Z+���$#-3��:VP�1��e����p��ؼ�j�ɹ��[?�]7|��kO�G��AqMOd�dh57b4*�I2J���>����<Įͳ�=�sӗ����T,C;�Y��J��pB��R�2Nr��w��'9*��u;�VU��,�b����[����_��?v1���/��s����7݂g=���W��٭h���Q�"m3�?{��>�q�>�t��s������K.C�9����7��g0���	�ic�Қ�5E��2>��A�&j��_��C{P���/an�"��~��ֿ(d�7?��8��]hGm��]���|�tӍx��~oz�_cq� j�Z�6��uo§>�y�&��A��K�?7\w5��18���\`���5��?�J}Sr|՚-9b3@1Av�`�� �W1"7l���� ��!->|׷p�Eg���y��/�Қִ:�t��E�X.��|����g?oy�[�`�E(^����شq3Z�SZ�ڜe��H=��/�?f�؉�����'cnF��Զ# ����*|��r]'2V�DO�k���o�͠ڌ�_X@�x'���g]�{��y0���w���e�k
��n���]���/�Kq������=�T��]BF�(ǵ�݋G���q�/�<���{ދl����3P��&�����2�t�B�qJc��`�D-�`���H�:6NGX�� �q��.�K���g>K������s�t�mk�c�y��/~��睳K���DTd�%w�w�Kv����ڨ0'��?�����w�̳��\�T�2^8s�8Y{�sU��`����LqcZ���b� ُ��{p��b3�G苇��g�� ���û���Ӵ%!��}"�u�%���M
�Y"m'�V�bW�$B� ��oԞbc�� �s����P�R"m{��;w�x�ەl�k����S���%�r�
�9R]"!�r4���B6w�zأ���R�h�����g?_��y����(GG[<����#��h��Zo�,��7ߌ��/ğ��r�v`������.�o�q0���t�����(���O�g9����z����V{	ƂR8LgZ�J��$b~�0zK��P�g��x��]�L�,݃�-m���5���bt�\������'�u�����u�1.����܅�/����w-�E��"]v)�Ze��{�ޡ6G/_@%l�ݚFczڪ�
�q0��p�j���ˑ��T�kR[(敫�����()z�ƬW�<q��m$�k�����eg�Ш��s�]���06��!�i�u��WkX��Y.���L��&��A4�����P������J�(B�6i[$V�	1E8�t�be��)�q��`�E���#�*c�cܒ�5�$�CZhWW�;�f��ލ����E�,uPW$�PqA���/�u�zl<m¦�(DX���%��7��s7����/x�s18�u"7�e�aϡ�\o�μ�B�$�+y�0D��-��}# >ec��?J\9��g�UD�'Y�Ѱ��[eV�(����]���n?�n�zK["?����^�R4ڄ���h��7�WA�A������mÇ�}�d]<���m��#��;�ȽL#I����\õ�f��1�qq�b�e�Ȫ'đq�S��e#
-'�&J�a˔aHvj��g:[����}�k_����0]5\�/|�x��_����y�FYO���r�x�uZַ{�yj�Fu�N�眿��G�i���_Q��T_��7�8W�����g���v�]=��>�1�3
�Z8���:��� @俉��N~��eiQ^����p|�<��/~/{�+133��7!�E����q;�6o¥��_��c登��Ba'N;k#��m��v��>�ױ��a|�S�ö��������e(d�J+�I��G�����`gxnu#�	5�Ɏ�e���v��ߋ��r4E��[/����ϨF)~��/Ŗٍ����1,�J���n�NO�׾�5ر�\����]���ۍ١�nD�~fozǻ�ܼw��JK�Ȼ�� ��Ѫ�(`�A/�k���S��GqD�y9&k��"�j�H�4���+�'#L�7`�����;���/���z�4ds��֔�]�y�]������w�@��x�k_���J\s�wp���ik�p�G��FP��W�Vi.��_F�ލC��8�ZX�%p��0�v{�5�������\�uō���1فn�������ô���Qco�/�S����'��ϿQ]w�q'.<{7�K�8�� z����`��ͨ�ut�4��׿	O��_��7ށ3�:��y�D��0}�#EK��Ae��ulk�9x�
�D�j�����<�1t�X�I�d\�h��H�6@��j��im
�� ������c�;����o��ضm�x5�Om�:��--���o{3�x�p�m7�='�h��7s@�t�{��:bx��<	�偅:w]k@� 'S�ud�+?��p��eK`t�߭�1Ҹ��a_Q/&C7_AI���`��D��k�����x�{��v��~���Yt�0�f��3ӱ����Y�{!n�I\ӊh��s�c��qסEl:�t����	P�q��%�fS6���qJc��H:�Ө����,����f0�]�<Ksg��o|O;7�3�M�v�=�ᰂf��5���-"B$.�]`j�N��&�/��K�}K=��y�r�M�v���cv�,���xg����5�c��5����\]j����w{#eW&U����&"1,j lv�y�
9fq���;��$^���?y�><�<l&���{R&�O~�����3p��O��܅�hl�s-q���s=�l٩�}ڋ�	z\���Z��4F9ֲ˖�/�-���,�k�Ĩl6�O�Z^�����*GKv���3 ���WP,����@ܞ��{2�a"����1�s0
U+hLoD� ��c|Э�9�S��uO�3������7p������3���r�lFD�򤯋��"dX��޲i��,�gsl>�ǔc���3v*��2 ��X�{ϋ�*
�6�y�<߄F}�V�Ȉ��+\�^�XԒ�+%��/��������ʗ}�(?o�]����0��ϗ=k�3����_�&����6�1d�;2�sH���/���*Xw�~o���=�����(ĳ47���DUm�D���"�۷Ga��6�R6��&H�@N�K���+b����#l��F0�˄�V�T��KCT�R萄�2�U��A�I�	p�zc��5A-٧�Ȗ�$�F�7��n_d�:��~��ZQa�t�K4�������>��(�jJ�C�"����/�ǣ�0bT: �щ�\���ص+��D���*��ـ��H���I�����7��P�C����C�za)[�g]`�r2�d60E2IZj(��J� M�תW:���"�-��"5Ɔ����x��/�Q:�S�a�G5R8�@��=T�M�1%�y6BK��c�F�#�r�Qd]�,C>��>Eg��{�������6�/�}�����/���G��Ncl�4/�**�S����ˏ��WǄ7b�µBy�	@�b��exGUyXe$�L���=Z��]���I�Mrg,.Á�M�،�j����>��.
C�ue��|��#�+]��/�4x��j\��u4�R<;;�o�TQ�Q�D�<*Z󡛉��T�+���Mm�X		Gz�Xo�E�J��.��A4k#�q�5�֌l�)�S��ƍ;Ā��� ��FT�<�ZA���9����)[i$���/D����&5rZ�w���]FH��MA*�̣��Z���r�X��?F-��lT��zA�ץ��/�m��a,�P�_�M�D&m�hRt��V�����J�ԇ�X_�Z�X���b�|bG��x��P�Ȇr��9��W�`�T�f�`�Ar�C�؆UӟS��)*������u
`_�YZɽ��ĕO���y�]����k��M�[�Z�i��}����l�09�Z=2$�9wؖuQY}�Y�c閁���$\��f��5��O�d�G���Z�v�7�'�v
�?&�X��A*$�_�y�AODbńp������O��Kx��_߱(�p�Q���(�INdc�yi�W��rqn�E-o��D�[�LP1Ru�Yjb.�t������h�4yds��q��ɳ��e���Q��_w��tu���������e�P��5]�7��H��}��nwZ6�A;��Lz)���פ1��8��l�-7�X����UQ�Ia |�%#��%��[W�����w�H�g�`<�q�Rڬ�R:M���ڥ0U��3���v�$�i��d	?w�&�ɯ���'��h;�R���1��͡��.��9�q(����兯����(0q�x�=r(�99Y��T��UqS�*C4�yZ�-ٳE����!R[��[ɺ����}���B��[�Tɠ0H;x�/�,^�a��)Ɲb�.����Rɳ��A)�(�(C�Q�VQ8�l^����pUk.�X�?���\��1�s n���&�ŗK���h�t�f�,D�<��Ύ�J�a�:���@��N!J0�D-)�6�f3E�S�c�&�&���Xψ���������í�G��ޗRO��yZ����EV
ő¡~N8QT8\,��OP���8(I�u.�ٝ��3���P��CA�-1[�㮽�`��I�N4�Q(dÑ�%y�G��h]�@,���᠇��ѣG�e��*�M�L�b^�h�t`�C��nCv�?p�_J8]�I��t3���[������(nc0�x�K��)W�=��Z�'�����:�R��>�w\�s�>�3-�� ���t���Ck�9��[ŧ�������.<ː�s{��+�5�������� �p���D ��j,
�+RGD��5r�O$Z�P�d,��TwǎJ�kj?w<���f�zL�<�w־�Ȁ���نc�{����9d��0�o�:���hk;��:��b#M�30X����VÊ�V�Xa���jk��П@���1+36�����%����-�Xh����;�/�e��j<��y*����V������?O��<q��cœ��P�{����=yc��f|��+��>�7��qC�,�s��H�i<��+����~���ص�¯�ʯ�[�:���:���'xȣ��o���n>�#�UG�%qp�R��e
c+K����Dt���Rz1ˇ�'z�/�Y�Jǡ����!F�mPJl�J�`k�����}����'��]g?Y��D���*�E1�?�����{j�i12E�U�8q��5���,��*�w/�Z�`V���3��*�ܳZ2eZ��D
��]���V6�S̠��`wP���	m����n���,�XJ��p�Vh��(����Đ.;���O:9�bY�O��E�#N�"#5�*t�����^���)��F��"�F�C�5�YNG.�T� �P������J�(,�c�M�h�,�6�l~c�3ч�">��(I��,O2��������'��ۂ�X��o������0l�m����>�)�+[��8<�(Z���D�b?Zn~Z
�k�5��Ȯ+���G�o&��z"͙��h�b����C�s�u�Fb\�
����a�3��^�
���U�ᘞ��+˘��h���G"�5��f;�h��"��s6��\r�$@�h
��	ϣ����A#Y�^QE^o����Bc+�7
����|lj?7P������rI��J��1*;`dń���+\6־8\�y�[G��X��,�l�Ao��O!���`>�����6o�푙�Iv҈gG��Q�1��i�dRb(��AilҖK��D�9��P�b����gU��A��F2Pn����#6��6G�B�8� Oא�;��zD@�%=s����I�D,�sLM70/�e�X�$�"+Q����Y=�0�a-?�+�0��ī��q^Tk
�dN`krĈ�=����r������13<'C�f$��10��^K�w^ V
���=nΘ)F���.f[[1�9�ƝmY��y�|řh��ܠ�	���{8e��^X��dt՚�x�J��h�.Fk*��j
ݩ"@���x�6�T#��Ē�n���.
c"U��r�.A@�������@c2�#@#�/i<�F�yU��pc��-��Cr�1
k������\�%�v���&�=��#�h]�jx^s1�I/UK"������N��W��c.��e@�9 5X'��2P//��ɀXbЮ֓=I->��AqQE�'��իG�⣂̧�2h����&����r��즙Y1X���(j	�"(��l�dCl�{ZG"�K�	H~+�H�ʦB��
Y�D��������r<��eh��6:8(�l��G���|OE4G*Z�뢥�X�B�#l ��h�	R��H�~i�dnR��ж��V�3�%�s
�h5��SLe��ĖA�u���S������A��?1w�e;����QrBC�U��P�ͽ>�M��t^��	XD��\jm�0�C���O�ǣq�mP)�l���"e�������/�,l�[@�w��[��/NS�4 	�>
۸u���Ƭ�:i�Ա����%��IҤU[�z8g�n짶Hz�Rk8,�̉�PC-�Q$�<�����F#Nb?��U�X�{���b�ʭ���"�Qè��+a!L3�>�шvz���4Y�$0�&�2�Yi�JA8�`L�Q^��`Иn4���c��˼b�Ǣ�xlя��v:4�������-[eJ��p��()�?�aV�G9��8v;��	�L�ٕIĞ^�����t|ظ6n�����&�3#~��{x �;{������b;��g<N̪ȃm9���t&R��&M��/ޥj�,��f�^�|g��.A��NG��^�W��"��QPs|�EC�Ӛ~��q0Wk�QUW�8�G��}Ypf+C��(�]�F�-gwU<�@Y���⎒��L�	<���(2�Qs��=�%hb��#t�J�͗�raA4r�UU�WmY*���2Cz$�`��N�}��jr� �p.��Z�X�����8�b�{�����"-���$�h��!��vY���g�� \��?��!�N�[��J��� �L=�Bŀ:p��Y��?�!N:��qAA���E^����YK;����h�m6�_{Z1�^��x �ZZ��6W�2n�bw$�(�X��RO��b�k�"U�Ĵ�@���2��j�mlajX�,(��|��.\��de���%�V�P�3���9-ǤQ���%�F]V�#s��+��$��0S�D��Ȇ����,Z�`h�%-i�V�e��nte��D��-��]&�LŒ�ԵK�=��@]�x�A\���fԛ��W��gd�]���_��p�E�;e��C䨠��` �;�VE\�,��~����@��ކ�:��@�SC������	Y���p��h�� %�!`�
�)E�i�x��³(�,F�h4@�M��G��b�*�R�T���a�̆y��)%	�k�.����}+SQT��)�I�+��"r�����aE(� �b�����Y���xW5�™,�-�}�E�GM������yn��p,�b`���2uG���W��r�����8~�B#��4���ҵ�g+�" ���S�x��A�!�Hu٣IA�h�*6EC��"Ҙ�H[	y�e��scW�cQ�����+�ȃb�?��NTXp��b�G7U�4�IHEJ㙂�x�ުB�����!zWd��"^����(�m퓖ss�V��v�5h��p�H�s<�X�P�8�VܒO.�R扆��}��v�s�X�	wR���,�#^���S-��E�D�]�㸳G�Q�jq99��yD/D�!�4*.���q	߉�J���>H�5��w�r��5��hFa�I,��,6����Q8�\���q�VBd��zRdU�x�$o+p��Oȭ6�xc��:L�h�Ck"�$�S���Ƹ�H;1�SӚ�]�,�f��)dؽW3�|e܁@e�\�(5Tb1[U��bYeq��xz�Z�X�`��!�������$��8�1x$0��դ�Bn�(pVK�\�x��ʻ.�'A��6�=��1���A���Z��x���Z u�:��w�`��f0i�p��5 �K0\�^�����9P}�P��-�;$�6��*v��OML$Z=�~W�c��g�f/aK!G![�@'���{-�	�P�6U��rn��e�B_�q��	j���y���P�3����(B���#1�#CS�C��e�X#�h�t���o\��>J9Z1Ĝ|@*�6�ۊ���-֥�����Eq}�u᫟�\;o#�~g���/��̣-F%#�*8bwt��҇?n�X]fkD�Ϝע�:X�9=����]�>T�9#�N��'�e6�����E�u)�U&��8Tۤ��^-p�-�a��Of��A���"�zMÓ���u��Q�4�џ��M[d�&��C��w��ϽL<��z�i�6��Gj^���1ƪ������%�F�g_��~!ww�Es�K�z'����-���i�]Pm�П����p�Tf�k0;��v��X���,1��-��>KZ���U�Yո`ʅ�X��銊�dK^���5[H[&&��>���_Ʌ���(�R:��}��m�g�]��x�����/GO�d��d�����~
ؾ��6�'��K_{�֩,f^�8���dԣ�j���[O�U/�/^�2�6�@D29�?x&�?�g?�J۩�2��^�y�Lm�Q����_�_��'��h�7 �4q˾%��Wc����jaO�
T�G��5l\�����$��8�A!gK3��M3�X��7����G\����Qk��n�����n�\�+)Vy��5�ח<�I�͙a϶
j��~��E3U#��̆vY�KC�h����2N
�KK���}䪲#1�2����U�`{b=w��k+�B��[� ���Ɠ�������2�F��%i���u�#IG�G���B{%7�S�SF���B%yr�ꮲl@ٖs4*U+$�5e�f����T}��j��e�㗭Ze\a�Q�߿ҋ��%�EVVÛ��f`!���ES��H��9Y�,;���^����=���.������o�#���^��X��_)����7Y��2u�NhT�L�z�/D�����Ci�<3�GPZ�����ל��u���MvT�n�����ǆ�ѝ�Ul�l�dM;�f:�sW�r���5 g���Z6.�U�f�#K��]��xմz�aC����Ov ��x�2f��X�i�/�հ鍜�}a�e�{�uZU^�Ҽ!ih�8��J�G����c��	�����۞�o��o�uzX�R���Fk��+n(0�pƑih{�=HU�+��`<��f�'�2��D��7�B��T�pe�h��,�dWOq�C[��zR�86��j3���� ϗ.zY����.>B4�qBϑGG��*6F��-X�6��\���3B�[Ȉ��s��pe+���ɱ_}G�T|qn)%��I�����-������Ɖ
�FQ�wN����윂�D���V�[�����١s�=_�ڞۄ�s�;�q'(:#V���?V�1֮[-Wb����2ʨZ���{��S�6%��O���y��-7��+��WV��<�Iן�5�IL���;78�����z��qn�iP��լ��<w6�� 'c-�k�v_OC3��3K#>aS���
˝T5���G��u^��aBV _�� ���|p�dJ�C��]c�T0�^�ޙ}s2�K�Ń��3�%�h[�}U�c#!M��B��%���᛺���6��u+�(�	'~V�U��:�*7���=6��;�jh�G��;\�N9�8�}���7��0���bh�Q���|��sN�K��h�u�����l%YTKX�HT���(mP�:��+��݊@�D,a�Yq��F�y�(5�9������w�E�(Z��X��aeO��S�XAUo��uP�;�2��Lk跢���-v�l��e��&4���U%�?Y����Di���r�Qq�,+��,D��!���(�4�oB�r��_�_N�Z~?�/�)U7�I8� ͦ������̿-�<�k�"�]�ܮrH�YK�c�M�����(�)���e�Ga�Y�G�]��I�`��W� ��}�}��4�c��љ�<�w%5�Cd��4�����u���5�m�w��ǳ�����}v�z;�[ Ѭ���q�A������w�,L7�ǐk-�Ά��X��_#��l�(�� ��2���Ώ������P+�+)F}DVMA�Z?����ֻ��*4��i�NT�-�����0���,/���|��~��ZB�G�ח��$'uKqƃL�I�-�rN��1��(��(1�n�[y�z*YD,��r��s~W��Qva�"��h�M�ǲ�w{,�>���Q&����O^��m`��ziM༇�S�*'WY��_23Fc�Mkڊo��U`F��ベ���a2V1Ũ�E;�wؔ��Ga��^�v�Fd�&IZÜO�<`�Yl�A�>&[���� �7����Jo�w��+>�[�N �w�&�<L��������`�s-��U��"i~��!����A.G��,!]Y��΋�}��w11Q�V,�.�(\s".�MD�-=���m��d��jv�{(�й��]t��}'&j��-1��Pv���sx��������!O�
:d#U���b^��ui2�]������%,����2L{U��b���N�aZI�f��o:�_N�������c��ba)JQ�aMI���LU��L6��}�6pE�>����T�0ꃳ*e�����KP��;�X�T�βD�<*a�4�=�������>&����W.�^�%[��ܡ�X�#�*b�,��M���Qf��>��Z�jb���F�{U��Rg��+��=:r�d̪��i�v���}�C���
��+Ǒq� [���̝�'
����U���51���`��2.)�[%���Z�2Y�`1+��P��x k7iCd���o��zݎvw3�Ċv&�<܏G��I�;-�W<�������pYH���1Zǆ+6�0��j�JcF����:D'�jMk+r�īh�^��(o��>ܰ%��z�ݥv������Z�����Im�ͱ�
.mj^����la��\���̚��H���Jh�~���
ƭ�c���G)�f3�1��%pY ��u%�WLElMd2���Z�]����N.�/�5�c�����B�b�l��zl�[��!q�f��'�Y����c��E5d�����HG�?ʞa����i��q?j�]E[x^���X_�f�z�5��|�++����ވ�Y���':�6F�6�[E��EI�(tP[��U�D�S�:�y��n1ºz��e�~��p��K+�L���fD?�J���,�8�N�;;�Z��5|
VY��&�J<�td�
dD���ŝ8��]폰�{���9>+�u��AY�V�W�� Ř���}z~����.0'%�sS5Z��Gꪎ�q��C-2He���E+Vo0ޥ�$�U1�3Pau��XSd+&���4�R��ͬ�5tF�.�b�Vv�6	��T�KSm�]��z\�'��h���h
�E���r�[\��v�-6�&������Mc>֠�Q��EaU�
o���g؊}&�}�7��M(��GG�E���{ޕ�-��mP����y��cj'EiN������a��I3$���@1��tǛ��D��(��'2�$����d�5��U��E�^֘fV��F(N�h0�`Ҩ?R�B��,�Б�Ԙ9ʴ���i��H�LB�S�90ΨA)l6g>�vߎUl�����(�x@D����x�q��H��^}�@��|h;�g��(�[-�T�`XYs��D�xP��U�6�ar���!�O<��� w�"�r4vY���uВ3�a��ݪ��X�����;�&�|�f�1�F�q�s�?�fg��.Y,O��X�^^�X-W��o!�~��J�ɝj�������"�(��v��������]���6��*e���H��]�j��)G
���h���:�*��l��#�0NZ�)n����qF}�"��^����C�*�o5��ׄ@xOfbh@,�O�4ǘm-p%y6Af��k����4L~c��d��Ǉ�K�s�����e]�0��m�L�c�*��c��ǸgF�r&��~��F%6W���^g��k���C��/G��/j�k�5���f�M��ڮ6�Ѱ�Q��B����jL�+rx��
i�Mi���Q�.�gv��|������k0����������Ñ�� s���Y�8@-D��i�X��*J<���:BWk�,k��S��f��G�w0]I13a�]�����Y��k����i[q޹�cv�F\�5���7@�kϾλ���۱Y�%�-Z�1-�G���Pm������hh�r��r��������bBN��x��L����Iy%��Yۨ�	�j��qе�Du�S0�D1ĭ�� RN�I2��3���(��.w�Ot�H%��Ii	�6M��W�;������x�_~����ٴ˱z�^��$���V|������֕"YS���	;/}8n;��-;��Qo�����8��4A�q�iC�D�f%,r�I|j��ʚ�0\�D�7J��v��s�@�F�4��¥;���M8`Ho4*�����KbC]�1�[-5�r1�'
UƑH[�p!�X�V��\s����ѻ��q՛��z�c�
䣞���Y?�0=;��z�x����o����}���O�7~�٧�;8�8m*�-�0�b�����oEy�c�T��Dl����}Ѯ#ͯ����.()���_~��#���O�R����@�*b-%?��Ǎoz�|K`7��JW���Ko�����0�˞�r,UN�(n:��,76�a�y �A(F�ᥡxm�%$�Z����8��}�U��]��k?��wnr���թ��:��=d`�������?�?�����Y��F�L,�50Ԟ��:��&a!������]/8\��ڒb��a|卯uu �6;�|n�1�����bg��KQ�r��-2�H�bB1��kk��,��+������`�\����L�A#Ws�+���D����ȣ~�"saU'��v��tw��O��M�۵ �#���,�1�%�R�0�Z�T0מF֛�L��x��G���6b\=� �c_�_f����8d�����W��w��k��U���/�����Tis�ץ+�TE���@0��s�ծNe왠$���&�Ɓ�:W�}�ӱ{Ǵ�0^D,,.��`��  �:�����u�=ޅ����	��,.��,?|N4����:K'�@!������p��	`dq1���dQt��+�VbɤV�"di��S�aK�ŗ?��x؏?��P!&Vl�),�D�q���B �@ql%��ۿ�CK	���7��]��,|/]W
�}0ֆjE)��������T�Dh5�sS���X�$Y��j�1e�]mn���-.��"���K���˰�T�⚆À� �z�D�S�������+�6���d��,ʩB �F���gl�o������ܪE���Q��~�z-���(&>���!	[M�6y����|�3��~�|�s��O�|/GufZ\�B��x��d"��`y����3���R(�>;�"��W,]$.8��LOOc~~KKK�29<6�Ɏ����D+�Sf;�V��/N s���U��"@�{�^9ƕ��*!�}���1ը���V���w��� 65]<�I5lV�bJ@���G�����Ǩ�V:Ǐ~�ݯ�E>�=�hO��ngQ+��j� u��V����	-�c�!����E*\Wq&4�Yg��Zd0�(���f�]���녣�U����r�\�;vh�Dwq���H�$n,�6���w�]�y�'#ɓc^��lLo����Gr�d�{�5x�c?������Kt��0(�������2~����J��Z͚�W�B1b����ݟ�'<����A��ʱب��*�m�~���qz�y
��%��Y�R����"�B,Sn�ZՐ�Xҹ�D]aR���͊��:�_cȍ�s��W��5>�G�+b�h�'�Q�gq������v��!� ��?"�LLg�~�C��O�5Hn�F4G�i#A>��X��s�A�f�������H�!���~�9x�[���={6�G��2��r�I,��]�ڡ�J�ȴ�g?�Y\��������fu�J!��ح2<��T;��q8��v� �4;3��
9 �L���©��&�����׆;7��׾r�^0���Ƨ��SM|e��(B��G~����\��wź�UMQ9�,��	��6Ÿ��E%GV��U(	��2ţ(�;wlBk�6��zl��n�� �S�����ᅿv\�(Z�%Gk�`��H��SSSG���V��^A��v�: �D�)=��� ���X6��Wr��䓟���k~w��\Th�E����Ck'�# }'ល��O�9S�����¡��е9NqL��ۉ�:���P9�+2*�+����_w��fkZ���x��Ql��b��9���}Pkl��%ફ�£x>�h�ǜMX~F���dn�U:-��^�?��G�B��)_S�щ��s����6X�B +z���y�,;�e	����O�����Xs�ꈰ4KW��qѹ���������%Í\� 1�Xͭu�.X�W��TN���@�	�C�4��G��hvW.�ԯ'FZET�pi �0v��c�_Lj�ȴ����~R��s�?|�׷	�]Y�����]�� ���I?j�8��5�4�fx!e%:��k�������>|<��'�����Õ�������*w��U����"Sm��Ts"��ߍϊP��L4|	��y0��6$*�&]Y�ǔ��=�d8�,C�h8���0N�/��ึ������K��+~�yY��cbpM�h-���ʮ�m��4���F��6+��:�����E[�k���J����1�!(W}]N�Ĵ�ߗ='r��a��@<��n�y6�]8&te�_�n}�(ߺg��-�5�����(��&�U-VV�z�&F{����J��v0��J�ܠ�*�ipj��q�rj�D�+
l��D����PR�zlGDLۂ~�ų�AO�\���Z���+_�v����U�A�3ϣ�+�׌�`��>�[vs%�!�[u�z��~������7��O�w�d��/���<���1�Q����W��f�b��.yG���u7`���jk���MOa�)Ζ&B�+yI�ڥ��k�7y�H"~O���q�Rڷ>C�B�;f��M����;��ٳA�c�Z�i�8Q��]GW�b���v]s�r�s�N÷��C�lQa�hvO�=i��U����%��佒��~����C�B����u���B"5oU/a�ؤ:@�Gx|�T큲L8X������_�7�.����遟�.�r��VL���V���Gj�uUz�
����V^�q�E[��I��k&�F	enS3�J�=����Z�kaLIf��W�����˗���<�"-qb������i�b260�7��e�T�r������k�ť�x(~'ݭ���G���K� ��?V��e�	Q���G#wK�1M4D��9����'��߷�B��/����ԅ�vaf�z��Ny�6��5�e��� �#rC�;���P�� 8v�C&<6nj^�a����q�RBS�#�P��Ʊv���Yl����/��.��C�-�}��a	rd�� %�*�rKN�
�:T���	��S���uo}����@�ܢF0��T�r��T�
7���Ϗ�j]t�3�D3�L��4�n5,?prV���=�N�3�\�	L��iL�X���`���5�̯}�B���i�a��(߻�?~���_���k��!q��(M��f�{Y>ծ��ط <�g��e1ІU_�k|%�Kp)J`�������4��zJ�{����	���7���"�G̘D5�S���D�&=Z�a�QK�ԕ�e��!��߲��������[���������]�e�Y�%-f��n�[��;$첋��Bޗd�v��T&���/�G�����d�ғN��=뻡l�R�"��|��/�%�_��(ƅ���:��`Y��XV��h���k5,f�i�$.�]q�Ȕ~���.6o9�����َ>�����=��.6������o�lR��_��P��U*H}dB�v��`�ⓞ�Bl}�Oc�3ppd�ܲ�D���(���D�f6nV���?Q�梫��̳X�!3�r<uʌ�
�̕GM,�����S99�yX�s ���.���������蒋A����L �/ڍ��QhB���EW��NV�yB�=�]NF�2�����T��E�lۿ����E����^�
��߾NT�����5厐P�C�^�2�z�"�*����"�k�	��?~����#��Jt��R[�PQU�м���G��J�<�����\��G/:y�*K	�(���,�3�0�w��OL��o�t�����b|�w��=J�F��4����"p@��2� d�l�$V	eg���S�5Е�Ui:ɚX�����¹|&(j��/gI��P� �Bԧ6���,pѣ�����7_������YNR�{hb�c1,k>#��g�Q��[�x՛ޅ���7�G��=�OCM�)�$�C�Pu��G��k�,��KAT-X3�P�@�GvnnN4ƒv���ڼĎi /�]�6
ׂ��\�(C�c��p?���v����+��
�R,�Z-h�hX�j-��<`����$b"PRa� �I�"Z�0S�bkD0Y�^���/�S|�u���7_���b�T!b�E��}>4�j��V�/�O^�B�����|����H��1�V����u�@���ص��%䑙"&W��sG:�l�����w{%��6�T�v�T�5V�?����S���:�#��*�\w��!;���Fy�l�CY�Ly���RO�>1���� �Zؤ���#�Fz4�!Y1��.ϡ�
Nc�1:�Q��Hda�"�ڎ��<�E������az7��m��������z��
�ۋ����%������`�9x�o���v��IQ��E"�X�A�K�lP���!�C8��*��`Q!�蛲��Fg]�����P���nʤ��\��{�Ur������Z��f�20��&� ϱ�aB;첱<)�	�յ�-TV�*'k�7.u�|F�?��~���)=;ϊ)<���ɉ�]��F0�"�T��dd�!�HH΅��`���~?�x�q6�x�ȿ�7�x6�����`�i�7ƕZQ,�o]{>��k�;��
8l��p�C�{S{5Y���w_c8�g%܂�Q�Z���"涊��xdvI���'ی�,q���B&�R�,,P�ƐH�]�j!�Ո(�#��ȵ8�e`l6��']��+��8�.�RXUKк�X�ьR���Ri�j��-�"gdC�}�mŰ����k탇(�G�4S�E�eYZ�f����[ο[K��;o����x�k� 3*������Q��坿o����z��6Av�p㐣�	�F�11���L�3�9��xt�8��!c4g��8A\ Q@Y�fiZ��n���������<��}�{o�UTwu���)�����}��>�������Y�S6�$��'7?�=[�Q��n<��@�V���[�K�#:�����X�.:��U��W��V��Z3]y�����r�)1L�}��F�y�ݻ��k���UW����/)x��d�u%�-�j2�8�/�����m|��FB�C��O���9'r+�Я��gj�;�뱃���	����b�1�������/����1�-��Y��Q���*�l<��߉���S����ִ�҅�ƙo�0���7/�Щf�hh�X�s� �tUL=�#D�n��C�
9@SعR�8eۖ�"�g+�
n����_Q��9����&6]'A�-i`�QIٜ�1�K VYr���L�1m�&Y����O�"�%Gp��,�
���|�T��b�`"<���B1�y��@|!�V��vӱ-����V򒁉 koK�MOs1e2�`GC����K��d�S-R���S�qj����s_KۏW���r��Z��o�a/6�� �<wi~'��71����<�M"��
�JϤ-=�>#�v׫"m�X���|7#Y N���,�(�\-}n���	�DcV�R�`�Lf-�r>5��٘E�O�3SYe�FE[�C~r`���,�?�h�\�˼2�fc��v�1e��z��(J�J�kk�P,Y~�,���
�;��{�4)��/�5��cU�2����b��yM�Z�G�{���C�X�Q7%�.������l��-C�kj�=�^�L-h�-�b�pS��4NҾ5���e^��⏃���1m�8�������tn�
�1�.?,(>�5�S�ȹ_�M`��g;yߴ������b����l
�1Q�߬%cA�e�kMy�Ai�vD&�cx�J��-Y�mtd�X"I�E���x9C���&Β�OC�g��
Lr�q��5�{�հ� bh~	5b�,����H����	Ѧ���b%�ܻm9_O���!d��@��Bƒ�J�f69Y��U�4�
�K$Mc�6-�+��s�֢�U��6���t}�7ѥ�S^�d�X�}�z�6`�َ�	L5yv������\�/;�b����-up��r3������	�Y���B*JS������#!MS?��%�Li:����3iS��&Qm�jV���B�3�vC��3JF�A�p�k�.���h�c�v�L�u��%�,�����T��!&@�31O�l;��a�)�.�>ĝ�:jrjU7��e�l���� 7���+��a���o�
8�*��9G�A�RR�����rt'J{���MN�5��d�#6�ݜ��\a�d�D,�oX��;&I���3g���|>Y ����b�R�W�ТN���|[A�V
d��V�Հ[�+���u�Z2�Cc��:-(�؆�^j�����P3ju7;��6�u��!�ԄWC3a7A���0y�s��	U�0�N2�EExZ�s�����v�VdbҮuqX�{E�|�oh ��CՕp�	&5Q�X��e�f~��U'��z���`
����C�,��g:� �5���{�&��Ս�5��&,bm�h��h%�*)lH߰r��]���\�G��y�ͭ.�\��:�x*�sZO��vsm�@�+j���� �3ϓ�|8�Ψ�E=Nlu��mi��,�ew�|Q����r�)�A�W���%	��+'���k�Y1���]��
=�]�MPP�2�'���H�$���Eiw�Ԃ>hT3	�e7Α]X~f"�f��R
;���H�K^`��.��EK�ƒo��d�99*f��
�Ŭd����&���S-~f��XJ��)�f���Z(����y�٘yNgi��&��{�\ܥ�%	'��_|����ر��^)h;�o�P ITS"�Q��Nd�+MA�X$���b�,xWI��]C&� ����6�����{p��g��֨��/U�5�s���3�����q�a �-v�)}c��5_S;#*�}^4aQi��鉐6Zu�Dk����h���B��<�>��M��T���+rltŪ1����QI@�YO�H�S�/yH�eX�wԖgU$�<��;������d־�\��W�c�J�N�&bKw#���^8�5XV��yY��� �cS��P.�B4B�1d�\�2�RK��I��GP7Mz;�#���G���xg��4���Y*:&�T�B��&})���,'�MY�xj�b����x�ٽ���T��^�Xhf��d磂h���aW��]��y�0��F�#��"�%����a��5Q�IꚲG򋤖��H�%	wD�1������W��b�T[y_"��Si��B���٢���!C��G�g���*ʎ���F�HSi�S���MZ>(����ڬ&_�\6�c֓�4�'GFsF�rX^'�$bW[����N�7�7}�أ�:T.�Y�5	.)��/��7ɸ/bkfy��!,V"ylcnF����kI��`;09n�r�����,(�ʂ��y4��-WV��/��r�䰜"ir`����,�.��9&�����Z_�h2L�6z�&�`��;��P����U1�`��VPk����#aH!''psr�+^ ���9���rbB7gw��U��;6�QW��ب��j��ۗy!CEu�T�33"�r֋�*��k��&����햇ju\ k���1�����/�!y��'�]��T�sZ]y���VQ��\��}�w=fL�[az9Vrh�Mc�%��ИhCu����(:��%���"��u?0AE�x&�M��=���:�
9N�{p��c8�����0|�i���-���<�\l}�)1	c�h�݁sљز�Q�|�|P	�e2j��a��2���� ���5�#��k
�a{W0E�1"��W���k�И�����ĝ�������Gy[f"�ΎB�w�F����ry�蔕(��("X�>���{��`���t��L�,)�;1ʲ�W!��Ƿ�<6!�{��?N<q��.��8�����W����/���-pE �����q�Y���'�C�<���"L�\ds8�2R?Y��XL]����"���)z=�eQ����L�8��g��W����gw��t
.�����(�[������_(��)yE=���k���k��O\��\v��j���D��t��Gb�Ƚ�2��;d�����k�;	����������F���������^�w��7��~��r�;X7���{���{p�+���W��ct����+�a�N��f�&Wk3�~�p��+RS�없Dc4�r���~u�����K��{o�[�r%���3����%B��޻Lͅ��!���YGs��5o&��o
�'��ʳOö;͙��a	#u��h�Q&�TZѶ��M�1ˡkhG�J�d��1���P|����ӂ��������o_{>���?Fm�p�ӣ�n�S!�>4����?˱*��=�c�����m?��-�&&�+�1�u~م�}Er��D[��;�߀��0���"�I�"��B��.������L�;��s��-�:�����!f��{�O�Dy���ˏ�	�굸�~w�8(J�!|����g&����v\��w���l�	ڙ¥g��~�;�\p��w��ߠ��l��s��1��k~�
����}��(.��;V1G���.$QgqGփ`��M�D��y�u�Ȅ5j5��qf�8|j��ȏ��^DZO<��%��wn����>Q��h$f��\��	/74�6[CT}�+���(&6���^3��*:/Ml+q�����σ(����+O��:'���~��9�:���ߎO|�2|��7�L5߸ �07ׄ@̱6u|��:�k�|�F\��Y�M}b�E�g���$��Π$�xσ��o��ٯ�ת�������w���;n=�Qǋ(�R4���U��tF'��\���rΠ�Bn�Q��:/�����]w����β���׏�=덣�W�O㸕�䬔�#��[�S<���8���_�"�H���-y�zm�6[*!����ΐ�jc�R0)�ֵ�v�Gan���D_�,�˱t��S��xIP�`���q�
�:���߉�U���Wn�����������D�4�z�E�4��T�ڢ��N�Pm�ͅI0I�&���#|5<�Z�Q����������.y5zH �h��a`�����ȕjJ�ҳYKIN�Ǟކ�_�U���7q�2fĢ��E^/i8N|�\���,����<�� ���y6�����j;vlǘ�m�=M4��q�ƺNǴ!�ã&�W^7gń��l����<*��J�*�OU�擺Y�p���73!]��O`V���Ę�B�%���7ނ�Gc���R�c����0Z^�����߻_���`ƟϠ]$O$�Q�+�=L�މ�+����4�W�*���FPA^ݖuuOn�!��\��a�9����w��:��ΚXh���v����ג�[y�Xe9L���E`b:��RQcIGb,�%Nn=��X���[(���"�ڻ�ֹ8�k�u�n��|5pꩯŽ��BvbGk'�]�m[6c�3L��p��ER��KLy��Zr���u�8�4tF?���X�UJ����b�ú��bӶ]芠޽���J���VKZ%����v��ǛE��
8&&�"���|^�g�h�����q�[~�ݹ˦��"u�%=6@��v~35������;��4�7=���j5yt��wc�Np�l-��gZTc���o^��7�{����X�Z0�Zq�H�\��xP_�Xr�Ĵ��m�,��a�7%�r<&f�f��L�?�p���l3�Yg�ؽ��!^�oz��}'`�ګ�G,�+.��>�"�>|9N���e�0GrX�k�i����Z�ZH��t�n	���؃�}�
��0�v�Jƕ>�NΥ�	f�9Y����u_��?��I&�g9�¹��A]>�����o�����;Q�2b�#u�G�֘�1+G�H\�T��b~7�|>��_·nK46N
��]�㲋�����n��j/��W��y�w��O\���x+yR4�tξw��\���%\�\�Șah
�֓��6BKH�J�,z�����|6?��y��V��A�����<��^��?݅��;kN�㺯��]�?
�z�L�|� �;�߅�b�TG&ЊM!�U��N
�ɍd�c|r~p�#��&�]y�&��]�ɗ��^�-�o����L 	J(M��O}�Q�Ys<vEں{�z�$������	<��^�i��V�1���em��h��h����Mw��-<���P[G�-�?���pʩ'�7 ��~��=�1���?�c�uڙ8���`/1oxRۓ�z~+J�1,�^X�8�Y)_�c�0�����J�7[������U�}���Ҡ
�6nA�H�}�I��ûerD]�{<Y�T&��z�V�{�"Z"��<}�����N�yL2-�X�t#Gf����t�FmǊC��ZA��06=�F�m���y��&�{�!�6b�����>�r�iN4LՕ'
0���P��N/��61���c��0��Ąn������ڔ7j��ʽtEM<�m/���S�L!V�	�� (O`J��]?} w���L;�ȊI89G�[���s�a�B�n��b���J=�.*�5��07�f�&�Lݣ�95I������SutR��YdS��Y���4�b�QlZy���8x�X]�ZH�E����f�V��� M�_!3�=�Ֆ�ntM9�b`�R����{O���k�e�6�aƕ��[BI*5yF�¸��W�8��mkg$Zn�$���wCK��_�Gb�n�BQ*�I6�6�r~(����n�����8>����2Bȸ���TC�j�m���fՙ,�/�P�%��[��$Yu_A$���j��9e5z��:���lƒ��<p0�O�g���fFj}v�����hn�>r�os:L�j ,�,#�VEw~���S7�8��s1XRijK�L��.��[(��+�6���8�9I��+Ô�P����@��*�дgBNfڇ�R*[�]	�ѫ+IM	�YN��k�H̸dȘD��A�f�w`��v;�?D&}/���6|�,1]1m+%��wuA�W��>��,:� �.�9r%���P��"*xn�/0ĲH�%�i����3YעB���1�"_Y/X�i-ñ���Nb�gW+�px4:ME:i��r�C�%�]�ˑR�g����4-k�|6���AH�� MFnv����L'1�_o5ܒ�0^��q�E�1̙��>����%�D X�����m,??���n�G1/��4�5��}�}���[��(�=���0��~ـ����I�Ք:h�<jXGܙ��_�N��=�S=6`cv�y>���{�s�[�����g�M���Y�L�C���Z�GuxT3��-:bAl�n4�I�T��w�ƈzi�� 2ZG�3FA�^]�����_Y#k_���Y��K��Bh�E%�d�%˲���~��k����U�@�ڲh�bT��G2�)CLb;�?��ɩŶ�,�~i<3V���|��	5�[�N��~��:�X <2��,\ʉ�x2��vD>�P�F<��M��^̳F��l�'X�7�XԀ�G��K��YMg��؆S3�dwT�t���|�������}��2{� ��^��J�wy�PALu&�v�Y��ǒ��,�a�t��J�����f�h��ҋ�9�\D3��i󖬒l@�M�`
۪UK����/�ݬ�Yi��l�T�~��lz��m:T�k5�,�\�[�[�i�X�	��y�ġD��L_��L&��TL��M��fǓ&A��ep=��\7�f��$j7�a�Sd�Q�PP�D$$E�m���C����󥏃���1�ť���c֏r"S�?���5�f[i�>;0˫c��E���O��n�8����3� K��h�2��Dq����[�J3h��.8Øb߮:�l����P��hE[�0Ɏ��T���5�A0�\�J~_Mc3����J*3�=����Ũ�v���Psj�\�T�Y'jj��tvvZ��e�Y�+�0$p��.c,�����݁ߘ���R�BFJ�M�S��I-m�vc��u��j�|l�8��i�]*U�7baP�n�,VÑ]W�(��:äh�h'�����I\[39�HLN��&GՋ\<ϵ)�L��h���	]�^�B�ߑ���g����#U$Z����=�1C��Sj�����g�7�I=F/����� s5us�����"�֎��쎒PkRY�C"�?��ۊ�]m�j&��x��<�Y�K�+:U���k�t��f�f��,C��5���c�%L�%���Tr�^ʤ�G'He����v��R{�� c#Qqj��z��w��ۨ�b�G�I7����`�E��8�'aI(�t�~�i����1��uy�jf�.���jO[f�����D�܍Z�wш�9����~Cch�]��fn�5�Pt�&�DU{����/�FzS�jo_�s�xz��tP��Ư�g�!���j��p��?�-O>e�J���e�%�ݘ�1��4�3�d���Z��\DzL2�~���$��a�Y\��s�n|�~�j�l��Ŗ���0��B�%�ϬtP�{te�eT^�bM(ܱS�����SN�\'���$J�1l+δۄ��4=]t���B��	�X�UC,&��f{�+VL`�ʕ(TC%Jcy`�e"������ڂ9���V�1��;�Be���W��>
f���n��L�g�Zt�E�C�d��I�Z�Ƥ��zH��q��VKwp�
�U{f"�l�TK��0u{�ڤ�1j��hʢT��-|25nd-�)��U��wH��1?0�5��G�O�n��<׀�N�!ɉ��P��R!w�[�$�J���!��APNv����Z�S��	v*��FC�ZM�����[��<l�!A�K#�9,<��A�M�7Z���o��p�f�W�>��
Z�϶��rrg ��)=�CH��}�J�{B��s��'iڗM�jm>�(�M��e掺I���	��YE���ؚ٬՞�<K|;}W׿�wA�"��Ts�m�=ǦO:�ݲ���B�S��jwǦ⩊�S� �-��p,ڎ`�PS���L*;�\Em}v,�r����N��_�l�Z� �g������ɤ�ϜI�`�g�zb,&�Ȗ���v���G2�ˬ�h@S��3<���1�*Y2S�Q�iE΀X��Ƭ�����hu{~�Á2<o!�J�@��]���=�6�<ƞɈlNbx*L�(GU)���Sx�hV��v_���a�}��n���ps�0K%����K�kL>�)2��*�%bIP�źP>V���׷�%��d�Y}��\���U.>���YI���j5EӸ�T�U�`9fU~��'8i��4ѡ5e��quc��D���$Y�Q��f����4�~^F=f�˘m� ��1�	���`Ǟ��9L�U�]M��,SW�)m`�bH�*�}z��2�s�d8����KQ|��U��٨��R�\*��@�VIg�"���)���xP&Z�`�I�Q�X޳���S�@��ݘ�������A��C�=�m:��i�����g]�f$ڔt�8gI�.�(a�gԣht���he(��j
z��,S����������ʨ'��MicS�d"Q���A1fيI�P��pkʱY��H�-dHk"�Qά���f�i�bF{e�:�b�ٽ����1��Z���O~.��mHfg�b��"[7c�.R4t�PvB�S���gFN,���4��FMP&�K
��{��4r�u��{�9�t�qfy}qT�gO�56|����~g>�g�����=���
��bQn�>�@�'�t�5�fo6��o�Y�)�\s�k�m�d ��G��f )`B���S���ȏ
���=�B��i��a"�@�0--w)IV�jg��0��3-4Km�je=B���d^[	Oש�B�u�NS�V��
Y]�$0�����ޖ����2�$0:r#�Ly��b�fy���p�H�e=�M��3t�Y� �D6Dq��
�m�HyRR�Fj�����ܘV�i�΁����P�ˏ��t�m	�����)���!i�l9H��OTS�-�Z����I���+5�:cΣ�.Q�����NK&�.�2��_��+�{�pjd��[��\�<fe#EE>��06���רFI��@vl��x~>�D }8�y>'���b�_������J_�fTE ���$,������Q]�mnik�x5�g�@ǩjL�����S�F�l�+j�԰�e~�����*�[Q���\D�*������{�pN�4�:ن<��X��.�U��@,'1��b�9%�˫А��jH�|�Y�c���g��� G��`��t3�4_�$�4�i�D3M�}%�=��E�@D�1fs�����	ztݢ��rSC���RfB�D d��_�
x�����j�tt�o��;��m,]o>6�GY����x,�NytT�挋5|m���pJU�Ϻ�cȻ��E�p�Eb%lD�Qv�f;%��2�8�o)��9���N�xEF6Mb:�XFY�܀����9;���Q��M8$J���&|��;�"��l�*�\���Z~�d��d�A���1�;����_�����j]�p.��e,'����Q��I�I���D)[)�4/�-:2�,��r�Y"V���7,s"�*�zu���� 8���u%{N�k�
�d��'M�O��f&����۠)Hb�VB�9�T�ihW�*h�A�(���ޥ֘�?���$�+0�6!/!���`w欦�65�ɓ�yyͼɵ�^(�/C*|Ij2�� d���u���NL��TK�r��Ӂl$�.�3���0f�%�R�JD�%���s0&���G`�,��؀%�z&3o#G�5�-�:(��+g��/+/k/�'�0ǡ(�f^�C����k�(w=8��7�'��Kר��-��p�Zu+k��t"s�U��O�AG@n>ߑ�5���"��vC��	��0A&(1�SqR�������f��O6�Y�T�+�u���ԛ@�SG�K����䞺ih�H�^W⩮�0W혓�(X�A���`�.8�RDCE6M�`�]�-^�G�rd:6�L�w�ɵ檓�I2_ej�2�s�r�5��h�S+�y*0C��ɤ���b��b��Uu�%a����[�=E�u�[�9����u c8j���cCs4���|�/��#�8$d�]4SB����=�;m�}B�{�N�i�`�+���Hh8��	4��8�<�иè�e�ш-���X7��	-'�̙�Yģ�ڋͳK��Ԉ�蘒��`Q�}���ibx�X	mG1	���E^o���3�Q�T:�}��"['��,�����Q�nhh��:�M�I@�fV�(��\��ȘoZ��(�{��q]ߓ#�����6�v����5�FNO(H����b���z"���Wa$ECО��B�]��X)��2�<�ג�9����O3�f7҉ɸS=]k"g�+M���?��S��(3a$Z����d�b����	f{�q'	�'uc�IO��H9@�U���J��.`d	�����O�V&b1@�s�`tc�\7�ϹCb�9i�T�Փ�CS�x�ߡh��Wn^�"Q��y?�Ė/jy�Q��p�-TGdG5v��D���f�i�b�;���9Vx�DF!���5NJDǸߍ��|�:��sI.g�.�0B��F��]Y�Ey�1�gŁ��j<�q��0����h��>�h̲mu�K�����{�%��A�a��e��1���T�݊�ĵj��YBN{'	،v� 	��ߗ�):�޿c��C���׼t^��r<G= ����~�|�=��m�[��"�yG�۠�.�Fԏga �!���W=��:k��� ��Ҵi�E�p.�̟x�BŐ��ۋ�ʊ������H� I㚝h�b#�^'�B��=O��@OuQҸ�=H��5�����������S�v����Ǣt
�>Wұ�fKE��g�G=���C��Tk0�<���v|�ǳ�Ug|��z�0�[q���\vT>�|Of�4~��|+V3��h1�Ӗ�Ԛ����
�o�ƻ7�MC�9\ks3N�&?��������a�El�LD����az�?�隴��/��;�FF�l6���O����?�p]o�k;w<�X�Vav��7O�����-��M���շ�cc��x�ٍ#pm���6�s�|�������_L��%�\	�\��_�η�������������߽`>Ƶ���^��7,w�,������۱�T������9�\p�,�а��r���߿�'����ј]h+���^�����6��f�v}����N��/�(�l�Y�c9��P�0�(��8��_��:Ђ�a�S]�k�A9�ꄫ
��rX��2/?����A��D�B�GqS����Ǳ��)�1Q��e�x��I	,B�l�Q����c�ޘ(V�rf7��/F6��wʬ���֬Amz�����n{E��n�y��W�57s<�q�K�D�^�Hշ��q�qL	F�T^YL;�3�U2����ɏ_��|w(_*�_��bg�b�8�4ʗ
y��d�/�(�cJ0:����8��b���0q\vC�>�sD�'�v$ʣ�>����e{�cJ0d��O��xK'�\�p�z��ue�JQ��'ը��7��q�	�<��4M�M0r�eJ���/����a��A��˭��֣z�k�����Gl$��KO�^�؟�`���8�#]47�aG{.�0KGq�ɘ7D�� ?�C�����R1����O?�`��w�r.�����V����hjO�G���ڗ��Xf�8��_�c �l� ;vY����L	�Qǔ`�_i����r^�c�1��U20����5�����܂1o-^��c�s}�Dq/}$Ird,|��_��1O0�Y��s]�h/����e�d`̋O,��V�����Q�,�bj�Ʋ�ǔ`d~Vl��5�?D�Aļ&��I��|�M������Q���.'���(��m3�	�V����jy�Ϝ#��.�qL	F�[fa��o��,H��lCCCڈ��l.[ȟ�����5���pS�Q(��Z�P4E�NҞ庶��z��Uv�zY��-��2��cC�,��]�V��Qǔ`\|�ş���V��eq��1{�r]���/���۷�#BY��7��n,���K�X���T�3r�8���6�o����q�eU���8Jc�ڵO�ǔ`d�h��c��W���3j�    IEND�B`�PK   ;j�X����7  �  /   images/2b66d102-ef9e-4dde-8ee7-817842500f7b.png�XwPS��� R���PBU�!��B	M@E)R tH�J�^�JGH�.ҋ�PD�@QJ	
�}��͛�����:{�{�:���={�8c]����dddtp=��YD��
p6z�d�>��zh226�s���v�^"������dTg	�E2�3v����3 �)������7?�s��ܒ�G��/�?�مg��EAFv�o�{�/�}yU��..��=��} �����ɋ	�F��>/��-+�>�1�Z�%��|�����p%��9�#|*xPݎC��S<�'���o�9�^>�W1L�Q3����.�Q��Օ_||�*~d �֋��'uy��j.��9Z�*� �u��+�>E�� �U�L�.5!>�n���f��f�q�7Q�>��-g�_�T,�X_k����>�:�c;����F+��g?���r�q�1�����Uʰ���r�S[0'H0]l��?�הۖrm��O�������98��W�8
�}�)��;C��r��3���&��?�.���d��ƛ�d��M��X�2U:B�72���/l�b��!�#8����G��d�{��x���m������#럀�(����ū�e��}��� }�g�
�B�!��R�����R��QD��z�_/�)��1@�2���X�L�d �IQ�l���Fb� ��yg�W�o��t�Cy =�(/O2I)IGP�yYr����?"yd�{n�y�kΊI���;���!����jx{����QB�
�����8/�<$���9_�B{���H��w���;�a���S����!EK��ű���"���l�4kf�Z����Y�5h[Y���z�_Q59:�eɔ��5
�Iu��qV}��Ԕ��� ����TH��.���F���b�	�mM@&�cA��	�)�����mگ��wD��M]�_����Z�)"�P��R3���Õ�m��~�y� ���,[=lo��� ��8,�Lć5��63�*(L|�H�	�A8h-����"Ҍ*{D��e`ß�Cy ��g\.�PK���$CX���U����a0|�.Ȣo����G��EE���Ϟ1�$��|�B�ܵ[֘hkת���(k
E=��/��-,�$bb�MLc�虅�/�6R=xW��4����ZЋ'R�Uf�8n$Ⲷ���5]P�I1ِݰ�C�d��{I��M�7��B�!�P%�A�ml�A��ƀ��$�R�zi�pT$5h��h�p�V+d��<�~`pn�Ȋ����	@7=*谭��x8-	�v�'4k�߲t�]�Eo��ʍ���\~5c�U��-�Y�Ԅ ���D���҇ӌT�L�%�I<�X�(�,v����Wn��L4����P69����'8�r�rI(�d���`�G0�G�14�k�:���
��$(�;���lEo�y�B��^z. Ul����i��n?	���L�{���S�1'�:����\ϴj����^P".�� �]�@�d����|�� [l�T;���|^^�+}T�{Y=мJ��x��]V=�IS��7D������o{_le�@x�0<<�e�R
@��Ʀ��I�Z��W4'Vc{Jq�Ukg��ʀ=?%e0W�-�TT=�	�!�fy{o�-+#*�S�OH�)� k�F�,ѽ3�L}k���n���G_�,}^]�Ԉ{|������yο-*7����U�j~�afh\��^"��h�!�`؟�l��?�g�MMc�|�S���X{7�E��!�����r�~��ۜa_�}�p��&��D��%q:��~Wh���05����v�7��Qskk�
Qf㦡!�og�%�Β��V��t� ^�kp���v73�E$��F-v^�.�*r��NbX�z���>r��y�5���+�9���9�֫Ƣ�z�x��]�@��E�]���z=�N����%~�.��"h)+�ѿ���k�7�W�u�����e�⹠�1�}�?��V�v�@g�Y�a������%���כZ���a{?pt�n�3�j2\>�e(oí��8�*��e��CU�sf&�����3�R�o�^=���ǡ�^1Q:V�n�z'B]�4"Z�\5�zH\ݭ�1�q\7�2�H�}������������O������a�	k��\�1������ȷ'<��S��VئҵJ���`��lu�f���tAK�a*d�$����f����V�8�zK֓�z�V_C��kj�g�^�l�A0e7��F�e(�͝�ga�5��i��ʘWk��zT0�MH�	p�۴�f�Fƭ�EFF�W�4�z7�P2[��`st�c��:S�@C$R|z��X��#OG^%�/)�vr��i�	>�v0ʓ}��S�U�+�Nf��V?���[�M�RG�;�]��m�mG������2��;��pk-ǳM>`���`'��X��wTtB���X�g�/�+�4��Ȓҋg�c�Yh���.��7Q�0?���U�S�zw9W��C%�6�u�mƵb�0�+Y����������
H�h2����*u���Y�>(iS�(�ɷ����4B��u�Z+��0�����t)� � ]�I�	KoL
�l�y����)���L�whm��<��-��>��=z�$��"[#b'��9!��r�������OO�h��u��vuᑑ~_��i�����D�~CNS�z�흟J؍�Pfa�~�ϊ�xUk�2�K�� K�U5�B5t�F��z�ќ�l�zO���w.�{�oj��1�xlb>3��b��F�4˸�i�D���k7��UT�X6=Dv�O�Z�2��LJ�94, n��P���L �}���mu�����d�o�K ��p�s+�`�z�gup��,ڒ�J����o�)��6��u��dw6��m
�gf?���o���<M7(p,�b7�碨��_��נ��{�)�d��2y��z�ɛ�-�2�1�g�72�"�r����k/��g���hA6�.*����T��IA{�P�4|>i���7=�%^��0d����J՞+����y�:j�I�h8w�OT�n���^�^N�s|\CZ�劻�Kp�zY�3Q�):��źC݁
��ƌ 42ji�*�}S�!�"����0V-ӧ;��e���:k����U�d�w��[\ȯ��dzzz�>���e������ Ґ#	�Z��N>�����R:C������@����ki�����e���j��1�F��\���?�J�<Q{�rO�����B�1^'m�����A�d�X)9qc��ai�w�j�gN�隄�>s
�\����24������5:��(Ǌ���d-�ޓ�=���rT�,@,d��FU��E!:S~���5|c^�-;-���:���X�)�4�M���*�0J4��n��Pa��o���\��g��ե+�z�[�)�o����Aw�f�KpK3���蘏�<���Fi���O����3�ҝp����,`-V��͊�5���EQ�n���y�!Rey)�ҵ���վ��9��j��*��v���j�Ǒ�����`���=�&��h����8��-b6m<�I��nq��9��Zb��B%��[��n^��l�%�W�۶��O�����)���pa����M\̞A_ix�쑋 џ���^�!��&''g!��x���">�V/���1�__��-H>���`l�;!}0\��Ee}ˋ�n�y��:f˻�j�)��� x5�K����u�pu�F*;p����%�@p���Hj�W�Q\����W=��������X�����Uݒ���J����G��ٮ��J��� ���DB�ʾ�����4ܡ/���%$s��5�N�fj�m��$�_RYu-�*3�gdd�J��l܋�fz��ʪ[��'d�U5;��td�_��?��ų��i4���� /5~��&b�.e�"r��R�2�Ƅ�A��FE]��%2δ����7+�,)�<��N���։]�ϯ3"�u�R��y�<����h���g��A�hr�ʡ�A�W9(�&D&��7���L�Z��$Ξ�o%C)�`0Sg��L��m�g��u�`W�ISc��W�|Lc4?!�4�ֶ�R��$U-=�N����g�r]�B��pq�ʒ�32d((0��B �{�,l%N���F��s�Cw����_G��^ʰW���ǜ������tsSl��͖�ҹ�q��W_=�[�	F<���N�5�Fc#�A:�J��ҩ�%HP_O_����X�����Ș�[&����y�n�-A��C����6���w�(y����N�a[�<i6��w(��q���Ige� l�4n���I���V�Phfӎ��8�tw*)�����Mӯ]y��Ap���*���#�������4��bq���snE��u	\�V�i�/PK   �f�X�zm�B	 �
 /   images/4b3ada2b-268c-4f4b-9789-7d2b3b5aac60.jpg��eT�_�6<�� ݌�4H7#(-�t# ��!!�
H�HKIw��C��3� <���/��y�}��g���u�s�}�^�_�� <SSRU`aaT��2�5 �ѣ�ƃ�<�'��88�xx��>%&{��������3Rr
JJJ"j*
2
J���`a?������ŧxJ���[��O�r�ݱ�X �H��I���@  ��	֣����>,hxx�����?�ڐ= ���YP�1�{K<
���'�
5=���6a+�|*jZ:��\�"�b��R��(*)�������[����wp���������9.�뷴��Y?
��KJ�~���7465�����B��Gff��`�K�ͭ�ݽ�?��g��K����� �X����"}���?^X���[@���,��L�=��9�P�
����|Vam���4��&;�?j�������#f����@���pxؤ �V�g'�gj�^8����@�y
�������9��H#��;�����\��8��8��C�.�!����FG��w�����$	p������Ł�-c��Ϝża3��¯��ߞ�D�܏�_U=��M:�ts�\s�_z�xm���?�!�%1�C�>r&܌�gvk�\������������ഭ�t�������E���Y����k��+⟙{�H5zYN��-ڮr� �\m��)����>x�?&��E��cw�!dY�����N���BF��n�� 1��knA�ӮJ&��G�;�tC�J���]�)�ƪ��W�m��#�0�k\����zq��ޛ'�?�2���W���~*j�(	�H�i����~.4�Z�R���1����[�V�s�[��C@��uCݏ��ψI&��=DM9�Kf=�����[@H��E[0&y�b�D�g�����m�1��l�n�Z/ϗ��X���z��:g���-g��Fsk�n��}p&ӳ��y26x�g�q���8�~�K��$��2�5�q0{�^�])(�P��Y��M�Jsu��<�
xP�|IX�3�{�)[��O��+(�o_̛y�I{�IS�^@��2�'�y�n���r�S=P�/�/&��$���M�����w���=��'�m��1pE����!B��� Ou�����v����_��R�W��B��(��53g}P(@fqz$������Av�+[�M$"L��~V!��|[�Τ� �,BkM��
h ?�;z�7�C^q:�6�7��ۢ��4P
�&{M�	~&�$v��'[9�;0�~綫�Ϛ� T��4�1��EU\f����&{��4�\ٍ�kE�Ru�������[`��{ AH�	G�����=��j��Dx��׮8Ȗx���a�RFx�_ﯿ�� �f<�k��a(��	��hya���j�G����d�.�l���ˤ�����=�K��eT�����B���= Z��E ,��G��Z�nd�a��R�$�S�ϙ�'n������� ��Eg_Rv���R��=���,���?h���t0zc�Yq�f�b~�(�]���7�7WػOI��._�O�/�p��r!t� ǎL 7����~]BB?{8	'T�eӐ�{����4k���xrs��'�Ofms�I��X����X������y�.R��|�	��)^%~�dv[}¾�M�_-Y�;ī�(�,_S���s�2dv��o>�JK'f�$���ROK
��Lb"|��pNeB5��q��)x���z�_�z½e�ݝ���B����x�^_M��d���=�o���I��A�l��IeF�N1�������]�/܂� �����l�ʞ�s�J<�t�G&Y�s`_�&ʼJg��ҁB��|��|[n�W,�{��^B�"� ���ܼW��}�[�9�#lw�|"O<0��M5U݉&Y:��M��CS$�&�}�Ҕ���,�gZN�㛫zqI�%��, ͳ{]1=��/�>�hS�J@���W���[o�㳊�<6�5v_^��6�P�m9�}kI��po�7WOw݇�w�+^l�6!�b�(��������c��o�����!�2ф2|���Z���'��a�T��x�U�*�>���"&��\��7����gM�'��f�����뉋�y�N��.�����+��)�c��t .4�EU:��S�\֕��ڞ�ƥ�z�f��l�ÂTQo���RR�Q��^���E�7�d9h�u^���ԉ#�Pn�,8I(�bX�C
tn�vv�d�.&�uԉ+= �k9�j�6�^�n���}7V��x��F�o�R���E�{3��s�@w�ƨ�&�ִ�����ᎌ��Hm�y1�yD���U>�[����Tb�v���G�r`X��̎Y��GɒP��C��$v4n��!�^oɪ!ո�l$v� !3AS5i�S3�����uP��C=Y�~z�5�$�'�JC1����×�,	+�!rG�J�$1�1�9i?�e
ы*�c)C�4i�)���s�ϣZ.B�O��sz%�I*��J�|��N�"7:�1u��J`>��'�u{�+�pӯ��/*Y6n�k.�J��:�@��<j�������T\ �=|�Ѩ��=����1I����|s[*H�mE#�t�^,��ͅ�|�u��c��g�k�?~�ݬ\B�KAN;��|��ՏW���������Hc��A�TE�'Eb�ݢ.)6?[k��p�9nWd�$C�\�-�����d�>�6�EÜ�o�XR��EZ_� �.2�r���sP��݊[��|�4��nV��@\*�Si���v���Q���vC4+Cx��я���u�d��Y�e�\ k���eXk�"1U���BhU��T���<P��ߒ���2-�]dڃ���@dKW��]n�-k�I�*��^)��
i�ĥ�~����(F���Ls0稪8	r��6�hT��o� 5-⥆�f��Q�>6A�x:=��n��������7Su%�U�n�r�	H��ZŐ��J�"�oYo�FJ�V')�:�E;J�Rν�^����`*���e�hX\}v;@R����M�Z�|Q>���=攼%ѳ��`v��9���*~�E��k�C� A@�VGl}�w^�٦h���֌��M�C��nI/�+�N�6�{} �6tx)�_F1xrp�D�ӏ.@u7  ���s2<N�q�Q������Ig�;YfLE��Vo�GxyO=�ny�r,]��.[	��s�̋t�E���߲r�G$��ȑU�q�j�R�\��vn�:�J9��B�:Z�2��Y���*�,�g�IЯ��%F�{�Ϊ������PR�1�<A�e��3-�_����6%����H5��.y�@@~,yd:[�ݫ����)�j�+�����I�N�+�Zd�D=6��h����A�c0/�3�ģN��c��R{��?��`�؅P����o=���py��O��dH/�;V|�t�"��IIT������~�n^��hkA!�l�Ѭ�0�T���̩�I�iY|�ϕ��wk��\ο��ual`�Vl���!/U�q"W���=�1�c����v5�����/�m����<��;aS�f��ڂϟ
���t\�L����1�}I�	�08;��й�RL]0��	�4.=�6<`b�hn[n�>�溑WHp��^-נ�D(.%��-Z0G{]؇� 9ƣ�;<���7z�D�Ѝc��CT+6�o���$E��^��Xk���<=H-�����k��s��	T����l����N���N�)�������4>�>б��1Sv_�����5(�P�5l���Q-`�淭*4�HH�0�l~7�c�4n���v*��mq�kʳ#�9���,Y(��������0&!<�+����<q�R"Y��?c��E'���^-;^w�N�﫣�_��G����~L�;�5ɥ�%x��N����s���Md�g�'4G+D��J�iL����ensIP`�xS��s����T�4���:��#��QS�c
l/]M��~(e����b��bǼT�w$$���D2A��ˡ��#)��&W����P��BC0;2r#&��������߱��&��]��;ȋj%�q��/1 ����5:�����m��I���}�����eH~v����#���O�x�O>����	�+D�s�u��w���,��Vp�L�#�L���V�ȕ9���+2�-O'�&cMo���>�7	�0E��R��P;xKU�.�#�N����q���á���j��tO%o�VD��IT<+��$z�׋\w4gꪫ�'�^[�FA�.��%ɰ�[	"���#D���U4�D�7A�����B���uZ^8e�����(.+����u���e�At�wӟ> T����N:
����.]���ͩ�<�^��}�N�,3��2=�����R�|�=JBTS5�;�=R�T*M���w)�����#i������R-��:�Z�k�3d�o:�*���#�"ݗ�s�4����B��$������ZE�D�սAei�t�JXD��<�a���c9C�T��#�|Z�-���T�v�5�)��ο�揢�eq�8��n)ş���^�ɕ�=�U���eʐ���z�qbAq_��&~܇�>A�_#Q�#�柱�a���*���| ˕��]�%�~�a&�yc���.rCB:��4'��~���a�v����<;���9�y�t�	F7v�޲-��NN�hn��{��x���I�2� �y��1ذqK������fs�I���Ob9���d��i�����#�Ms^Q+'����w~TV?��,�i���$�K\-'�~d���_ګ��_����8	}~Pg~�I���o�t�>�r��"2�ȗ��A;����<�� ;�/Uo�z=��E��*9�;�vW�Gkx^�6	�	���R݃w��t���r��:+^�f�x�W�̌^v���'Kk���:-�҇�L_��L�e�����N8���sU�����I�+A,7Uq��w�Dq�m��A��k�H��HjVBu�}�t�OP@�'^p�^�2F�6;{+�󹬃5��P��Kb,��Að|�_�E�	Ϡ���SBd���rd�W	^x�5D�M[`�%Ԉ��h�&VF�~�:g��@����@���CPI��2)?��E�N��R4�������1�4�MxhԈ�W��:�OS����DA�\%bR�d�q�a�![|8*��49�U� �h�y�&8N���cm�Ay�)l�N�m��fΊd�D����[�IkN��y�S<��l����1��<Cf��m�FU`���%b�<?�|J�^A"D��5�l|�P���~��HK[F�rŤ���c-�}[��Z�R�J{���6�Ar��� ��<4�[(
�f^lb�Q|y7ׇ��Vә���qE�9��&S�m�nxzL�6�O,�;ڒ���$�;���s�(8�LG�����y�/���o"~u��(�,!�~6��`�/7!�l��5�?���@��u�o�Tj��H��[x[�I���6�%y?'*9Mg�>z�,���U��դ�^F�{$G��K�A'���c���\��+�w��\J�aX��I>r��7?^ٴ/h����s�.p���-�@��WG�I �����UUNv�Z�q �ޓ�;]��������y����Md�:�2'�8���֗� xj߰�S�F�|��WP��O����^Ш���r�{��#3�e+s��������ϛ��M��Fp��PR��?�+ib�Ǌ�z	&AU��$�ޚjbZ|�gO�'cW��Z`	�c���+[rA/�޸>�q�Ψ��q��;ʐ$9�4]�Rbr� '��C{�o���x ��m!�?㫟���O7q�͚k~:������îac̯5���,�
�������)�~��މJK�v�~We�sd�oéh	�e��1�r���M�E�S���qD���J��fm�=�C����:2Q׋{�ڈ�6�f h��7 p���Ĭo����|�QV����I;�\o-Ʋ#��*�8<L�	�������c'[���&�n��tLG���X2�E��`]�{ �`jQ!oֱ����G��Z�ߍ�������a�O�zN�b`�9hB:q'����{�p����l���4?3kٟ�۾vh��1e�f���m����Tٯ�S�����{齲/�Zr)��s�F
M��2w�a����̈�����K�|�T�������j��Q7!��#N�(�Q_L|��FxD���:
��r���4�R�(cT��S?��0���:'/���� �19��o;�ʤ�U�َ0���cF<IƱM�nţ.L����D�ww�4�a�� kwi?:	T�S�$l�i���˘|x��֨��tC%����ǲω�Z]Aj;����Nx��R�d"k[�����*�HU�y���	�W�#�\�TȪk5"_d{���:s�vƗ�T��X�GV�q���z��[������+%�==��M}L,�uJ]�u��'�-v��Lf��B:��k�i�ӼAQhvLEE�{�ge����͇�?[��
E�~<V�X�ŝ} !jD��	-�=����Z���H$m��~2,�<��γ8g-!Ψ��!�d��d``z����̧݁��}X'�]�l9�w�M:LH��m�׹g�{ �x5�#�IJ�/��~s��񒉥��1!0Snf���	S��������p>��5X`�K�[��2������M	΍/���;ȩ�z�N9��b�#�Ir5m�\���Ul����pH��iP���^����b]�zԂF�d��� h�_�x����Nbi�iux�q���(��Q���;�_/��d����|�P����$5����K�%	mqip����4X��3�fG�x�i+,���':���}M��f�~<һ�3����OKJ��הuR3�W�qJ�Dͤ�0*oU���� �Vy��Fzb��ߺ�\��Q5߸u��d���)NG�Ԍ:p�h�ֶ�he����i}�}B�v��jQ�D��#Y�o�=��+�WB���v���#�;����N� �+��W0���f�T�g	��"�t+|�0�^�U�{��FZ^��cW��9�%�<ɲ��W�n��@a�t�W�q7R�H�µ���D��nj���N���Ƶ����YhS��5z�V��X"��;ڧ��-�eż�7l����v�b��xA(͆�{�
������R-��FVG��?(�Z���m���ja}lV?j{�S������Af2K�G�o�$�P�����3�D{�O������wu�q�zgto�u���|�K+��D<�m.��rO'��A�)X����s�u}a��Y���g�i��噎R���x��Y&�ܹt�rP����,����8Qe��RM�M|C�@���D� G9��jo�?��oh*�}�,\e�GV·�)Mt�AU�^�蘾):&������yЌR21���3�՟�v��s/]��ӡl\��z�u�WU�A5�Q��"̓��sY���H�I#��G�$S���y�z�:�OL�Ƥ����o����=��k�C'�ӂr��;�x2'q.N�<X.�S��d��L�LU�ӱ�5��l���Yǁʅ� T9��x���\��Xj��)�������{@�S�
U|yl�A���'x�� m���r��!�ҟ�;���0�^����������HZ����,7���]���J;7ԧ�f:�|��+0���웯k��[p)t�)��J(����7�x&p[��<�;�Y��!����� [N_�����ÈOA�I�$��\������(����a�~W���q;��`��Ͽ����C8N>�Bc �m���!��>�?w㔧��	R��PI��_��͵��-Ci���an��GW8�!7M'!��[~'��Qr�Kb��J��H����Kz�������s x��ش��Uz���'���� gAtA�b2���46o*A��k�zW ���Y�k�ק�TA1ň�7��z�m*��m܊{7.l����Ǒ�FeAD����#�o�7D|Y^e�v�u�ƛ������L���R���A�	��Ո�+�|�0ɕ�F�`�{ !�K�fzn�S���D�a �JrK0���^2��vF��a|E0�'_3��[��Q����+�>�x)�1X���ܬ&�(�oD�)#�HM+&v�S��Q�xzY ��L���	�Kr�>E��𹗜�n:��`sp���\�-F��x^*ҫ�q��B�uk�_����)kc�l�L
��IW���B��p6=��{��ۯ.
6B.�h�>�\��S�˪����wk{� '�J�1�"�m��-Y7�:I���#e>n�N�I��2w�YX�%/�[��;�ҕ�얹\~�U���+������Hq56<���h�b�����Cv��5$k�J@��ii�A�uы��*n�t��Y�|U���g�\,�~8�PQG8F�PSG��MW稵��r�S�
SA6Ѝ�+�c�'z�D�Nx\�8�=ӟ�l�TxM�j�S�&S�{}�H��#|�����GF�֍�F��}Vd�^�į��)@%n�풟��:�
�q��I�寝v9�?\��{��wx>޾6�e��`�Jy)��K��F���V���8,@�����=�rӮ�z)FL�z��C�y�@�E��K�O�<[ҥ�������.t�>n>��i?X	Y�&���u?Z���ύ�O~F';ϱ$�N�E/V������t,���?��#i���d�������J��-����GF��N꯶�'��z�ee��W�ד�Y�_��GϤy�pD�)�
�.�o�~�Мj��[@h�r:� �i�`�	�����^6�5��7�����v�LP�&-=�L_�
!�G�5v��G颣"�R>�@-�&:�G�2 Kn8��5�ti���$�
�]�0��,Cݐ?�k넊Ќ��L�)��ޡ�3?2�egU�����s�ʞΥ��}Gͤ��_�L�k���������P�סq�C��7�JiJ����q�J�����鮶��+�
�Ly����]�ꥐ�L߈"� �q�2��,v/��%���h����2�®���zL,�*[���2��?N��$&�q��ܒ%����_)�z��jQ�38�G*��m�Wnb�,�5]:��4�1k
�$J�x��nD��(�؄xhʣT��kI?U�?�vMb3|�ȁ��q����������ft��7G��5-��
e��=�#���1*��$J+{��XN��}�l��1q;`	P%�3褣�y^�j:j���9y����Pb#B�k��}��{����M�8ԥW�nk}����DǕ��"�7�w0?�!V9�Z5�1.�A���)���GׅQY�M8���°&�Ȗ.աAH�eCr3En����΃s�e"i&�j"�X���v������}��϶��w�4_z�K�5���,��2�#z<�e���t�}�.9P�Q�҆?���z�9�E�v��N�uj�����л��/�#���D�y�Sgo06ڮ/]�{�P��.ap�75}99��p�A����ȋ�5ʌ�E˭\q�g�S�ľe�0VZ�]���sC0�tWmu~�_�a�<�ǌD�C�7��&"ҋ�w��J���bw<����ȓTv������Q��c�V��h;��	ϋ��&��_-$��>�B}~��'����4�����m����%.%ZP�@����8"���#֤�O+�}E�uЊy���I�|?g��$_��G��	T�w�_����\�㦟�v��W	���a�x6�x�+ޣټy�o�S���,������p1>�2X�F�pA��ɘ���v��9�f�''2���F�J��Z(�⮞c�¨��Mꞩm�s�]z��e���������`|��[c�o��N<�D0֧@	ֳ�����Y�ՁN��N3o�[4B�J�5Y-���q;�E�G�r G+���,�Q*���� ����8J���lH�9(�W�� zu��J�f��6JN���z�=4�qȨȁ��'���2RuU~RS�b��4����\�HO��vM�i��	(��I2X�����#��RgU-�����K��Ҽ��*?�~¸�H�� ύj���Y�o�pDɯG,�О$�琛P�2qm��Ci�8�V�� �8|9�Pƚ�8�2�A��Bן��/T�k��[�?�z�����͐�-�p�~�����4ԡ�0�+��Ҫ��W`��*�U�Յc��Z� kEy�P�ޚaLQ���'q��v6X�P'�q�3-kt7+k(I策oB�������^YRB�kL�(�+a�K�tz�vI�x5H��˯�t���ݲ�����`�&�C9��A��u�ǘQ;m�����8b��.�~�Ĥ�)I�炤�֢��>�a����Z���P�ǻ�o�ͣ�����(e��v��23%Q�nؤ����SwV=Y�k�������MF�'����>�ϪIs�,!�������Ss��l����߁���f��|_| H����V;����`Ȍd��U�I�U���S� '1��E^!tU���w�䤎�kL8�M��q�I)c�~�T�i�Oy6읭-(�Y�Q�ψ��p?�`�����C߈Q�B��_W���uk�Pn��w��&���\�&C���S���郚C������db�d�[�^W��_p$�FR�e�|�(7��
B>h��M��絠%�\�k-X�ׁ�f�Mk;8鲯s*��`GO�x,t�#3�^�����ߜ(+�+56$i���n�R��dV��*�4,|�ڿCI��k�����d��.�o��/w��o�>�e1�S�"�gK+���?��e�����s쌻��=Pݸ�P:^�P\zҜ�k�Y�D�$��>��Eߖ�ոˌ&����hh�-�L0���uG�[/8����|YO=ȭ��ĬP0�����ۢZ�G$L͗%4�SI�"�����ח��ѧ� a��`�G�`��m��t��~W1��>�X�]�|�H�>�Ey��]d�R:� ?uIݬj��m/aY��~"i��Tw:�����*i3)�4>}%�i*<�	p��ݒaķ$V�^��a�?	�CFI�~���ҜW
eCG��B~�Gk��v��	�>"�8Y�[ǡ�7��A.N���b��)��͟ñT�oEim�����"d5�y�/_y�ggɶI\s��\�gu;e�������RW����){��Y��$.��������VF=E��k[7鯕3��]Sv����J����f��P��	zz;v�e�������L#Wv�����Ɓy*�|g�`˹��.��Y ��E|�˺����)�QNX�� ������#��6�L�����lг�ּ22^��'�_in�5�x�T��ġ:Y����z�\�I,�Ҁ�Ilg�)�b��2�"��3-�f01&x�|gi�qZީP8[$�͡$��U�{��Z|�p\�ґ�[�4Z`�8��q����8Z��:�u�|�F�>G^�Ui(�8�}R	�V���-6�R�T9a�g͝��4]	]�ç�����X�-�� ��G�⍡s�6�λ����5EQ)�kn� n�W��p�$�x\���HH8�D�K�Cu,��P�5:(4!ܿ6(G����t�!Nt#e���6��6�Ě�.�!u<C�IghX%�9��[��M�q���"$��,2�����2�~�E?"F�[r������(I�f�يB+O|#I�ىu�<{X�����rO��Ҡ�?��'
F~��ߪ��#�8����󇻱NV�R��Gxc,.�X�pT��ϴ�uQ��<m�Gih΀,_!�l�T�f���C�3�}s&�ǳ �5w�p���)�2�>�>�~˶�ۥ.�!d�<�V�.�`�y����T}~�on�����Nok��P�ot�4܊9&�F��. "6kj<NoC#CxP;�\#v��ȟ�dm�ʹ��o�b������h�֬�9�e��z>�40r��Qb��+���w�*�w�����3���Jn�u;�!ԇ�����xQ gHӁ�[��N1��֚�;(nǙ������a��2Ĳ� rλy�t���'�V1C�ˬ�Q)hP��t.R
�i3�;� �Z5��Qҁ>�c1��`@�1�:IFQf���/����3���a��l%�3�t�<r޷�);��C�?~����y�L~���J��$��M�B���S���=��	+�+;
ŝ���"�+������4
�����x\khWB��:��f.�0�޾��34ߟ �M�CF��h���
�Kk�y���䕻�u����bД��s�|M�'|j�n�e�1aҜ��x��ZGd]���:�8���bs�������^��2E,�0
1f}R�?m1b/�~�y�s£z#�Z�����M�O���uB�KQ��u��P�M��<�ϒ�(�[[���u������^B��n�k�fI�uF�Zс3�}�C}��Xו|�}�6U�%�W�9$0���������7d>Z�a4����E�G�$�<+�"�?����drD�ѬB�
�g��N!����⌍�D����v9F{����UMY�U�G<�`ە�:���/%Lk)�&ٲ5�\�����]�^�K���B$yMH#�a���>���qW����b �I$����8����]�5�z�� L,��`7h�v�(�e�M�g�Sί�Lۇ)L�V:p���R���)҈��)���_�_��v�;�m�Ɠ9�5��̏����Ƣ(���Ƅ^�~�7("Y��J�xg� [ 9����h_1�{���S��272+H�t>R���i���f���C)����FT�ކS�֪��No�q��B�2����y%��y�'뵡���cݱ�2!GL�C�	��{�;U���׸������j���}���!Շn���q�S���SQ��	DX������z����·o=�>�ᝪL�J-�<����l�:�lM�8�x�v��
P�ڷZ�P�����P1Os�6[T�eb�mi-�d�M����g��|cP҆�%���/�v�$I�`��#�M����������t�=}�Ae��m�z�	��J�����z*Y�*1��WY�{�  �\N3���@��7'��!i$F��(��si����_���v��+ #I<Nt�X�xb^�&��s1��6�&Y��tfn��cT��Y&@�u�M��� (�٧��v���F�l�˚�4�4V�(.�r���`�p�k�⒑=Je�i��y�9�i[{�*�k��A�;�]�P`��E�,�*�ް}�?���O}5+���&n��Cɉ#V�T���=�Ol�V�#�r �ѻ��Qy���%���*���	�o�gk��L`�B��,�̇�={	Umjz,0Ъrd�mmz�=��AnH�����K!��l��1p�R�[�OF���o�ħ?�v�k[�#H��k�a�m�V�d�/��E�����q	 ��d��u(�K,���Qn8s$D���2��V�*��N~�i�d����x
cP��8��[��m�q��ǸpM`�E�)�6�L9�U�?s5�U���	Q��ۂ�]�`_5_�k�/��v3o��e��e�H�$k<yB.�X~X�'������:��Bw�����y��	�U��-g��iƱ��z�J����Fc(q׆�Rm���Ħ
�	g�.ٴ ���J� �_����9�8O�.��EE&�����kN�����E��*����d���m[C�Q�Hζ67B��*b�`�f��qd2_���P�4ƌ�hG��6�gkH���]�JQ`3��������fU_YRx�Yxm\���:i�iT�8��622PB/J<�B!
w'KUl�jCg���WΡ��>p�y������bVG��f�%Nz�do���0�c)X���H0���O(���.�_�}���xw�Ti��-'b��������3�TN�.����d[��]h�
��=���T�Y۸��ɻX2��ҵ��$9@}��T�V�}�_�� >�e����q����r� ��.b�M}��myOZW�C��ݢ�.�4�#e��w���{Z��&�/p�	L���˚��0s:�j��J4I�p�T�~%�i��"C��7%_��[���*h"q2�@>d�ޑ���E�WH�I~y����/ �u}D�Ks����E��@�W􉪶��/���ݞ�~CN���XHB���4��8x��&�sȞ��^�[hغ5��@�����4�Ȍh��4����^tTq.i����b%m��Ȥr ���� yB�)U�#ݗ�em�e��tZ��Ֆ��l0i�7&�<���֣�y�irIvD�}6��F�z��ɉ7� �#[~��Ml�G[�6����g�֩�;4.�n�� O���> �dt��g#��Ln.k���E2�>V�B;�TO|�������a�S��u�т�_��ky,˩��vי�J,{׮��*G��8c�%Bw�l�ݚ�=���A�NN���/O�:�Qy�Y�$�k�4�g'2��M\�7KK�4W5����0E��k�V%O�?���\aKk����ٔ�����Z;l��X8��?n��h���nY��U3�RR�F�l�ՠDu,�&߆����+��O�rg�$3�s�ƛ���~��N��<�^�k�ˋ�L@t���ޗ���"V*ӝ��ټ�D�Z$�������I�ڥ^�M�R�A�$�E������+�1Gg2��A~B���3�_l~�|�8���̖�����y �G�:�̊?}T���"��n><�z�G�x;�o���҇�jgh�%�H�}��Ve��i�ͣg���66�ղ����[�d*���A��j�:e��ظ�^���UØ�eV֊\�8�(����P��Ly�.���|���ȓ��?�.D�[Y¼��C�4���>ٱ?� ���*ŉW��=�9�ݿ(寄+�����w�קR��d�?������E���b���JMG�SF��ڣ�����yԯ�Q�k��Ed(}��f��n8g�61������]=���Z�lg#L�|*T�ҕޱ�*L�8K6懲�f`@�?���4�}#��6l��7c�%���z��=���2�B�8�k�rB8{�0�兛���	b���!�=oe����lB���~\ecu�j��l�/�u�#:
C_��� ��#�W�>�r��b#i9���w9g�~��h�6
���|��Eѿ�A���Q��F�R.'u�[�,�kXμ�˛`�m(P�D#xB꠰��Eޡ ���2.���TQ>���d������ 􋼔�U)���)��Ǚ�u@<�>qR>(��wML�#��06�W��*�#4�+*�C�̦ty� m��= 1-B��t�B}�Q����5��
�#6��Q�ELa�D��x��\*��G
c�>���c&��^��9��H�!R6�2�iuh/�^���{�F���<�p� ~p���۝����ʥ\ò$�q.X����6 _u���)���˔��=�E�G*;H�>�������aH���T4/����7�����D/}2!�oJ�%`!x\�Vn�_���1��ƪ>}�*���!�����R����Zd��^�� ����o����V͉~j3���>�!�!<{�`)�G�Q"M�҉��"�&%ɟ�6ߔ�Sڒ�'j;�:�оZѕ��y��D�5��N�x���T���Y�'xJ��6�]��k5%Dp�v�Vx(TQ<���􀔉^��T��"�QN!�?\&B�tWe����F��#^h`��������ȵ��r�Q-F�dW6�u¯Q�!����m�t0B]��ɀ)(�<��},���p:q�I'Sf0ؿ�E!G��[-��hK�R'N>�H�'RNgPd��=o�,�� ���C��]D�w��dmn�϶���$˙���h�~�lU�:���ܟ�)��qT�yA�x{��G&{tFi�[Q<#���d�=~j�HΟ�>;��Di ��J	ܛWiXpn�@h�����=G���n�u��$�%��T���,^�T�q�mxR���R��ĤU�0���Q%Լ�jm��hl�`ך��9õU:���O�x0����]e��,0֢�5w�*)&)��v�E�~"�J["����:����nX�)��H7��)P�=���&o��ӀEOR��������#�W���.h2��U��Sc� �U����ٴ�)���?`��= ��p���I��ȋ�՘�S�i>��n�aܕe�o���9�̌UB���z�M�o��F@?�v�a-t�v��(U����}ϓ(4���ByN�?!�%N��5�Ȋ��� �����k�*/$&Y��5l���O>E��|���a@���3��jB4EV�v����߿�~kǤ���we;���^�6��9�\�v� x�})��Կ��tUk�3���f�X^�M�Pvʌ�����'9����?��ޥ�����=ԩt����bxJ�;{�l�9���Kw�0<1��,[q��ܒ~_osU�Aٓ����)l~��SE�~%xgĳ|@��a�L�M�wv�D�Ȣ6�Ibcܪ���nxɯ���k|N�>���Q�_k����Wbd)� �G���k�X�'���t���~2G��>'�t;Y$�#�{�\���f|�s>J�G�������t�񶫡7�䄞D,s} %s�ǽ}��ut����ƒ������ ���g�R��=WO�q��<��ہsnNJ���� �}��Oh�<;����.l���<�u$ma��1_��)T�q��8�,�l�O0�F�߼�w�A'�S�zv�g�^kc�KDU�U�ЉNHp�����Jv��Xa�bI2?�}=>$�J����:~�U��Ga�ji��K;�ƫ�J�_�>���q&��g�L��� 栽���Z9n���"Q��޼���=?ᖗ��7��ά#�C��<d���j���6�qVp����˩J�Wf���_I���j���+җ�ׁ�ƷW� �n��.n5[���Ԑ���+���ӟZ�_M��B/{9
����>�(�@�)��~��kJ d�t�?�|��F�\�AX	Uf�0	<A��
��N���U�g��~ �;�#XW�>s<�}NA��~�($��á����{zz����𮠨5h !�A$k�B0J�˹��"����0��UA�ti��nt�*��r,Q�����5t��+�y8<��J)�C�~ў ��XkM�;�]�� �u�����kd��o�}"I.3����GB�#?S\=��Zjy��Y`�����'�$�=p@�+�n#�^�$��V���F&8C�.z��>���YPɰ�ջ����&q�"�+��,&{��j�����n�ٿ�:��].��[��gJ��nVgv����В?���-B���z#A�q�o㙽���Z�𾖾'�&�u�g�2,k�B�zg�y�m(�(�Z��r�'9��}��4���S�-%����t$<�f�K�/Ϊ̣<4hk��՟Qa3*�FƉ���ި�4����F�gv8
*y�e�S���1��q����u��
	�)4�R��W�����������W��T02�v�p:O�i���W�E��1��zp���N��e	M��\�u-[�F�#����۱�x�x�N?Ȯ����}�V̎21�u�W�k^-��������]�/"0�w�XuY��Y��;Nsӷ��K�JU�nQ�x��݉�&\>�Uhی�<Q���!ij�7�>�,��<��Mr��/t�� �t���Lw��|q���JQ�V#�~�.�+�&��I��w�0�ńmcx�]�-aQw�GkOC�>&^�᥸�.t+��$����Kjpx�i�:F�tm�ci={WL� ��ʛ�ðkr1���D��;AϞIY3����^C��pͻ�'#�u�+׾"|L������[}c/s�T��������6��8c�� �gk�"�th� x�#PP��q��x�㗏<U�i����_ب�$[ca�F?ɭ)�
���wૺ��g��l|K����MwR��������E��Ӳ��8!�l��yG����o�>!�ď#�>F��_�Ă@�ll�pA�^17��E�L�Z~��-c����:��1�ƺ����W���W�n`V̨�HO�c�#9?���6�OW�J���\���>5�|I{�p%���˓%�1�JpT���ֽ��� �Y�|`��q�iZ��D���2���G����������0Ы4{�y7e�ۑ�^��O�k�����M�H���dY#hw1��cUQ�=	�ާ(˚QC�j�)>���O���"������b�a��g��g+�cv���|{�s�x3᭞��x�����8��K�$�<�/ }x�]��/j���c�jR|ְ�Rysʀ������=�����m�|���_>�n��|�%A(�+��>��K�G�,=9%t|�o�|I�f�ӭW����g�$`^d��&vnnq�=�Y���-�Xx�-A"k���P`�����
pzwϥh�N����k6{I!�.4��6��ՙ&��r�p��W�.�>���@�,���l�16�w�Iq'�$���8�f��}+o�ӹ��*bv�~\x����Z'�<M�Ƴ��2�&�!�ݗp!q���1޲��⮛��/EԼuy�aH�RB�C��r�ǞO=+o�tY'�S�+x��M�n7[+H��2# ���� �Z����o�Kk.���'�� ��T�Ͻee�;������ƥ�~�Sxf��WZ�ŧ�%����������|���EƝ�?�v�OV�W�+����c޻�ن�uڊ�q͡}Ra�.]0���׎9������`b���&�Qs��O"�qN1��S��K�-��|�&�(n�}�� <t����l�,�]�l1�A�qު��ǂ�f�4�xL��&�T���с��k�S�t'P�6O�����m�F�J�8�NI��FWg�9շ�����мh�Z��5ݶ5�+�<6�⫟�׭�fY;)��A���y"�-�Č9'֓��q�ҫ���y��V�>�I/���3����3���T����l��y�?�X^J�$pi���/e%���ͦ��w������ J�7ċЧ�`�����X�B���Uy!]�4��N���5���v��
q����q�Q�H�3���7�J�q��T.�	Ppz��ʚ����C'4�}�I[�����4��o�/�H<�~i\�;��c<�k��xK^��M�x�E��uH�g�����7�8#�}G�����^�+���i$��ՀA�9N8�� ��9�����I[��UFOI��|�_ֽ�*�?X�?�E�߂?<}�k¾
���7{F/�mKǹN�:�߳���Mr*O�>"MB�K��r�l�d~u�w��q��ؾ<��g|��*kאE*B�hl��m��I�<c�l���G�� ��1�ό<sk��O���D�ґ2)�vm�� �͏��c�[�?�t�ռM��{D��wV�"L���O`q��QvH��p�z{C_�߳�_�О����B���ltd���~�Keno��a�H ��~ii�$�7U9U%����x�=� Jhd�t $�8��i�y7��>���~�z}
�2c�D�e��H^2�^�.���H�f�[۰ǖϒ�`�~F�����z#G����� �k��o�b�;Ф��\�P	f��h㍢�' ��q��s��+�ox9��/��7I�ǁm���`r�^�G�����W$��Sj�wef�@8�B���twrC�mRpJp0:t5���XB։��5��dQ�>\�9P7|�>n9�����q�<����kOC�/58-�V8�Q���FnN}q�}*���G�y6�;�`��4j��ݖ��d�m����"���?O�X����-�43`}�6�?�\f�5�ص�Q��o.��<���ڜk�#Y!Q���$w�7h�G��U���[�@3Ӟ��FJ[���$��/!����dt�1�x��gi����)`��V�آ9ݴc}/�$��y��Z�M1���̒=�._z�jʤ�#�R���j�!�櫣�VR���@�c�& ��	�W-l�y���P���G���~ �x�C:�������������;a3��8�+��?e�W�� [�W�|�0�Kua<�e�gz+&���Z�$���B�*����3s���~T�� q�qڻ�x</,�7��M̐��u�?RYmne'�lR��4{A�T��Ӭ|��`�&yb�*%� ����;����u��5�l8}��� 
��!��i	�$rR���Z��߅z~��%��+>C��D1�Q?�zc��YN���ӚkJ��nX?�^�{�?�-ucs��ޤ�3�L&�#_�����aާ�>|2��Ut=Z{}1�
���a�g`��G��N�#QŴ QAR��y� <T_iM���k���^���6�|����;#� �~�
�:7����J�
|�΍y4s���6�j���)��޹��3ɚ`ǧN�� ��4ʣ8��ѣ�[�Ԥ�mA��X��Č��m�ԩ���ib�{�_��#[���<�d��m�)�q����̒F�h�  �@^zƽ�� �-7�4}����7q�<���1pb�o^z��|)��u��� �,��J�Γ�˦&��[�"[�����HJ�'��S&��ʵ�i"�w1�� ��{÷���R���ppq���������?�k&���~�����$�Ӧ���]�+n�s�۞y�t� ��v1O�o�.�,v�XS�X�\\%��m_6Q:��� 0,���d�+<��q�^�H�px� �Ts27�g��i:V��MB�@����<��MxNБ�ߵ��9� �qX��R0rw��Q��~q�~���8c��Nl['~�AN�+�l�2�X�m����V�a
�c��1��/�S���t�nfFbs����pApل��:�C$)�8��.��85jݖi����ܣN�M�K�l��%����i������\(�a��{cңX�ӽ�{YFY�/�Ҥ܍�Lq±�O���2� �+ۊV�fs�8�42����ɥ[Yv�����`C'e� �,x��aU#��6�c��j�4d���ƕ��[]���?욍{��x�Z0A�y�&��u��*��e�����㹦2țVO���J�F�@�3�Xs[��s⯋$���5�[�i���S��,�(��@_C�g��1<q��h�v��ש��H�G��G��%��17����F������f�v���A״Ҷ~1���Y�Pc�<����;1t<ŦSg�� {���~��k�M�O�4�i��,�;bl�@=�F�����)�����˝+ůt3�M��~]�m!�?/�ֽI�^��}"�E�.�w�kV��lo�I �r0x$sָ��w>g>Nxow���o�F����ۑ�T��*{��_x#\:��纺�pZ;,HҨ���x� ���PiQ[�x��o��p��G��Z��[K�/̏��,�W���yRNPP��#�pXʸi)S��Y�� ��uf�a��	��DXL�o�9#����� �+�����6�MX�9�ʊ�;���^9�j>1��N��چ��%y=����l�>��o����]: Gt� �|�L�-���O�\Y���`�Q�?i����M7����w�]͔)�w`*��r���4��/<E�5�z�����6$g�|�q隭��1��ma#��ǻٱ�}i�-�K�R���pQ�
�0�>ʌ��g��Vw>������S79o���J���cҾ|��3� 
�|���I��_A��޾�2n)���}04�E 9��=���Lө�ҁ=��?/����O�^�;_�\1&zc_]�>R=��5��P��s�����XW�>s<��9�5H>�(�!9�Oj�V��i��G�� /oγ��_�L��mu��f� �B�8�ׇ��G�~��X/�]/�/M�m. �m�����A�]v��xw�֓[%Ĳ�cs>Y�#�=q�=��s���g�7؍9fP:�W�����v��9�.[deہ�~U�֭^O��[�ʧ*��3����w�h���^����ߚ�&��G�C��O�==Ʊn/�"�kqk�_sTx�\�#���=랤�Ge�[qN�F�k��]Dr��mex���x~�E�F߄#o5V%_�iֺm���_\5���ܢo11;�)���aU�I3O��.�-x�--e���0d���^�A��u����m.�����ck����$W��&��x>�O
Yx�R�w��J�H��$��$d0�❭|9�/��S\��w��c+>ۻ2�L���+�S��v~ǕaiV®H���K��� �(�=����F� ⪗�)?���$����Y�� �Wɐ��w ��#ќ��7h��^����{�b]�.��@�d�c�>�[�J輾� d��
|9hʈ��]M��~n���O���c&���}��{ɪ�3{*),߀��|��/��Y�/�tj{���׉I C��p����ǦxgE��5(�L��!��)G��"q�d�:��y��	�=��>:�O� ď�ڶ�m�}�j-ezC��Z�o$��]��-�֒�|y�$'C�h���?�/�|����^��g�k����*�����z�^8�_�Z�֧$��k��b{��@�>��j)�ڷ�_W����>�վ!|8������7��K_o,{����{f�m/�W�.>*iN�/�o�H.���m�B��ēԞ��|��uu
���ï��?�Z����9
���7.� �=����J�Hʦ�#�t�>���ec��߇�Zi--��ҏ�̊@I9��W{�ZC#��U�ݹ�^��I��^�����E���i�t�m_�L~��]��瓚��c~9�IB�pۡ�Y���Z#y��*�,�.�>o\��W�~�מ"�{�_ ji��i&�����Yz��.CpF2p0}�Š�A4s��\:����+�_�{^��_	�L�Eˮ��q�~vvex�t�%RVg�|P�����'�X�|�}�֫n/4�2[��NN텗 �6OZ���/x��Qh�Ǆ-o�M4�n�2y�2N����B�u���z�_��#� ��g���{��gx����|E��i����ڵ�m���'����1]�I+�H�P����Gκm�ޣuy-��t�(����{�w��Y�}O�u=VmE{��1�ycF��k��1F{e����[Ś�<��u+��yq��r��jΆ�kgx���C�NI-�듏Nݫ�xʼ�[=,��=��-�=���c�{�|'�(�FY{K��B:(��{}j]�ĺN���O����l�^鲤r�6�H���f�;�_������~O���l�WwG��y ����_۟����G��|���^�<U7y�{��i8�*�� ��|Y��?��6��}C¶�F{d�K9"�@�H�$�+��/x�-7�9�C �;����ߟ�����<H�|��T��$�N��|��;�|a�j�^�V�k�+��bl��8�"�9��>e��V�aNWw6�g?��ig���ɸ�;U�8H���v���-��M�-��o�t��bvn�i1�A����D�Əi��B�.4=^Gf{X.Q�̤4[�ç^A��ľ���.��xm�?a�C�yD�0�I��o^G ���ש��L(K��Ϣ~2�Q>�B�I��ue$b�	6��m�g�g�Ď��(�$�)ʹ����#��Z�m����D��>�ykm�-ĳ9�P 9�V�l�~��s�۲Y�ły�� s���^�z,��Æ�Zr�Fv��x�$,�*u��QI�w�쓓׎�=�Mu|��'���WD?(>���
r�<n����q�L�֗�'o��µ��MM��Ci���w?ʩ\���~�ˌs��Mc#I �U�n�/�ÚH��۷�S�H�)��}R�u.����V��G����|Mo��(�!����V� �Co+*Ƞ}�-O�Ȥ����ea�r�`Un��{��I� 1�O�k�I����'Y|"�����h�r�:��ŭ��o�"�޹��۞��s�8� ��~��H��k�CQ����qpm�qwu��'� �^[�Yx��sqqiqqe�� �����2 ���=�'��z���d�?�um��t�4腭�_i־]�D�]�0+��$�W|�l�ϸ�M҂�բ/� �H>i��|	y�_P��T��ye�=�2B�B�8b0wl~�3�7�?�Q?���!��!�W�]OÁ�%�����8^X�#d�a���9�k�3�67Z���-�d�������FV\zq�^���q��_G�x�:��I�+�Т���!$ڠw�`��+�6�1<E� :�m��?�V����UǅuO����B�$�m�fT9g�>��9��U��HL�����`���~�k�'�a�K~�?��/�wF��t��Smc��FDp���v=���)O�D�I�`	's�>+�VlG3��?���vQ�!�~I�潣�������O�:?�t��i�lma���ftW+��B�s��<W�~�߳����۟J�_�;I�.N���mo ��,Ī>*�8��C�.��]�2�3]x����>��߾博(�[�rOȹ�#�X�j_<]��7:n�d�.-$�J�����
� �#�f�i���־��ᶶ��͝����J��͑�Vo-��*� �A����/ُ�o�]������4p��I�HVTM�ѫ,q����������<��ݕ��oh��-���^�m��p����rp�־���	��K���k=�	��y+&A���{s�ڹ�~Ⱦ6��� kς����OԴ�_WhcԴ��\&Y*����1�}s�r=_O���x?N�u�X/�.-�-�ӕ�1����`rrX��D���	3�<k��Y���C�Y���.�n�'���dl".�3אk�.�����c�ᛩ��a[ɔ�r�1c�G^��x�ľ���X������_[]2M>�N��h_y{r�<ͣ#�1ϥ� �@���o>��k:։gy�7�{�@�806>SÌ�`��)FV�~G���6~4Ȃ'���nfk���^};w���_��}�w7�5�4�CK��R�-6Wy���j�VQ���}%�_��m;�^
Ԭ�f�]ci5��j�r�^k���e��pEw_���&�� ݾ��Ծ�4�F����i�< ������*���˱�S��$�XEpA��Uy�7N*9|We�>ebp@�8�=s�W)k�X�[s���}��I>�!T�j��1IS����=�5��jJ?d��3�������Υ`�m��<(�Av �lޏ�9$��<W��D��?f�g�i:v�4��p�v�|�b�!l�s�<�o�x��mu����쥱��VC=��HT:��ʡBg�O��������Xm�M+�\WfY!���ۭ�FĸEIprX�����:��΄ݶ>���u�>��'дmZ�e�/��y�y�8�c��u<�s_�K�A�]_xR���J���#q!q��T~�����5Ƶ�x�<�권�\K�<�S����^��˦�~�Q��4�,�WkuR8�>���;[s&uk�KbR%N�D/ ���\�Iu�iHRٞ6`VI-�Ě���$�L�ʰ� �z{�Z�$��Y��l�A���u�&ܚ��- {F�T���t~.�/�T[IVNJ*��W1o
M���
�m��~��Y���-���퓎{��=��s�(e�Y%�了x ���`x�OY<Ԏc
ŀ���z�?4ik�_(����}� ��H��>f?J �a�-&���Tpe@�02>��Z��Ŗ�+� ��c���}z����-λ���"��8���Ô�������f���i_�mF�������ݧO%X��G=~����oڣ�u����C��b�]A�Xlt7B��*ҁ�6<�p	�|��KĐ���5���ƑB���  �=Mv���~<�m��k�� ��}�E>����XG6�4cx->��8c�1��~x�}X��}�����_��<�|:���x���αb������ϴ��q�[�}=���.t[������B���=[�򠴒#�"y28�3ʀ���y�<4_�>"�}��~!��/�ǈd�-B	_M�8ʬ�o�2 a�� ەO}��2|{��j�:7��vi㷗P����{#0�3+s���{�)���\>$�[Kk�mL�<	�������H�X��3��(��8��?Ni���X񴷡/"�UT0�����6�{��!X23�k��~ʠcn�_�[�UrY�g�� ���|}�_�S���i�Z�yw��#��0�3���5z��	��]u	`�����V
�Ks7������[�z���=�d�sGj��e�)0�m�U'i�:�_;|;׵mgP���3\O�#��Fy �A'Ҿ�,�%�;)X�1x� �F�\�'�+�g��<[���M�ˑ��5� �`�K�A���#9�d��yB�Ȥ��ٖ�l�v>����������?ξ��uE�S���_�pV��L�7
�Q��Pv��3c��U�� ���8��~�W���e��b�D���7�g'�WԮ.l�k��yvlIJ����� S���ݹNN��	��BO�G�^>w�$F�m��7y|t��� ��?\9m{�JT��_�7]��uw�i�q��,~F��0q�ye�*���[����?���z������ �쟋8�<(p3� �� ����� ��������J����~�nng���F��?1��G潀�x�/���o񩿶5�����Im*�z? ���� ���*��})��k�}=��s8|}ݠy���^���o��8��]x����ge"�qs$q����1d�85�_��E'�&��v��u5D�`E81�˸�u�}�[R��������:��m����7�)��y�#M('9�'h]Þ+�3<�����wg�`�K�r�I�3�><��d�5��Im��Rk"$�)�H��k��aI9� �1�?x����#��� ��MN/#>��Ɗ�`2��~Vv*~�����O���_ k�8����E����Vm- ���S+;�!�U�99'�SK�}��>��ŏ����im�P�+�đ��0@��l�'���yN�U��!d_��i#T��~�%��N�g��H��y���`_��~-���}�ϥ]=ރ�[��lgS�r	�3�=�����? �ٟ�-�� ���sR��~٣Ãŝ�Vd�h_��ߠ���6��������c�%�:B���a���z�y&��`rr��;��6���7#X�o��a���f3HIf�n (��\DzǇ5�u���kf�=�w�x�;�s�6�ʸ�f� �r���2��7ːK���;��F���t�x� 6�,3�X�1E��l޻�����놓;�����'vq��Z�o����a�_�\�c�d����:�� �åz� ���� �^,�4��t:2۸�"^>�1ہ�_ix���-y|9�/�2)��a���7��U?q����"��#�<mm���?S���ۭY�ƶ�;� ����CA�o�8-��P�H��?x1�_�~��g��t_��9�ɯ!EN�g�K���l��|m��%�P@���� ��-�+h�yb�O�����ѿ�#���?۵����R�\G&Kt��J�eh�T��{{��)u9���G���,��s���Ư��-� �n˗k.@+��z_Q� �L>�n�G�5������<t���t5�a*�Y��bm��dTʞ���0�m�L�?a���~�K��ԦB`��3�k��{q_/izǉ�tp�H�K3<��lh�=����|b��_�W�Pj��������g����`�4!�t}8��W+���W����f�k��0��!v���s��P�+�/�\ծWa�֧R5Q/b9>������ j���j��a	�u�����|a�V���?����|G���y���<wT
n�-Y"_���X6yS�� ��WVa��� hV_���'y�~����㬴���.��W1�}�ŗ^�'�5�|9�A���3��W+�����$m&s�z�?DuOk�<�Va��U��֐��t�d/���iCv+��q����ss7q��Y��ԖsY�9We=��7vs�2�z���g)i�QI�s"=BD�͡I,�1I�L301���C��;9$E}��z�-Ԍc��k���~4h͎>��}�W���\�`=z�ߕ|�p�\%f��g
%<<���
��q�.�e#�3�_22��7\Z�/�k����7k.��}C��1���c8���8��*��1�P/��[�hΗ�*���[1��8���~���Y_��f��f�K��I�����Y�hˑbqOE�>�V�Ta�#��>� �Z�׍�c$�\��b�^�������}qe��Em�Z3�3��$g�_ԵH��vi���o�M�� O�I�H2�@�j�q8��*���h����9$�[�V>�ք�-��#�v��>Î+��~�p���Vň��JH��]���m
���K��|�\7u��S�����5�F4^����>����W>���h�i�c{5�1A"[K������ �Nț.6� ���� ѵU��,��)?Ҕ\��W=��cZ�3����_�#�յ��T�K���]̖k�gw�\G�4+�k�Ha�����]�a��^zW����[[�Y��ZV�W��F��f���FU���*�q�I�@Ni^۞?6������,X�������H�3E��)��gۊ�i�L6��94|J�涶��H ��Y|˧`p:�Zts�<��9�v��E6��P��O�\l5%%qc�m��`��:S.
��qn��V%��#u!����S�a=�pOaD�Z	�K&:i������q�5�����A?u����T�Q����T\�v*�ď�_��L{&<A��X\Yx�B��-��,�����dc5OI�g���4��mn�O����S����;�B飺UB�fc��p¦��Ǻ&UR�|�� 9�cRTU�����ڴڅ�8�=�iwqA�n�*�G�W'�2q�}��+,�7Γ�u7,��1U t�8���>	�������H�6�5���U���9�pj����/�>�/�;_h���̢�Oi��ʫ����NO#�}%dyRg�4�xז���۬�w�~��R����i�m�� c��� 8�� ����~,��S{V�=��+rݙ���c1ۭmY\$�~r9~ʭ�q��u�u�P��b��h��+�*Y��u����%ǩ�Tmi0� ׭+����Gl՝࡭�v���8�G�D�ZM��H&&c��<��ڥ�|�	9 p���F�X�l_ޢ���d�h׾��~����:�O-[R�R���E,&Bp��#��s[>� �g�2�&���C��6V�_ES��Upk�=7������� �SI�e���E��AR��8��4�ۏ���o,S�A��@�O"$f��-pJ�Y�䶧W�c�xѾy�����9X�D
�,q����ЋdgVt gq#������S���OZʚ��ƫ,�4�M�1���X>,��4�ǘ N�}k���Q�ٔ�>�>������Ь9_�Y�=�Ϗ���筯�4�8,�9=��?Z���m��؟����3�\n+�)���姐4�>����AZ�̡���x�o?����t]E_I፴���*.عu�`�"�T��|4���5�2�p���,��G��6���5{�-��$���2�[,Q`���g �',G�^O���$��aAǷ��Vo��\�#��1����v��+�����)�����@�Q*��(wv;��׊���ů�uV��@{�x���KAt!F#��1>��׾�Z��ϑ�# �۟�S՘J���-�~g�0��rs�����j{��3�޽���?�4Q��ir��>hƓ-�_)���l���;�7�����=cP�<K&�n-n5	-t��I���:em����+�u�����1�/���/��4�
X���Y߳I0���g?7Z��+�]���G'��s��v�F����M�u�2-�UdXp�e��qW%{�^���џ�C�]������\�º�k:N�yh�O���[�X�GFv�Z�<u�|x����7Ëh:=��6�nb��Z@e�D�P�
 9��M}Ce�&���� T����Ϙ��q�h�+ȗ�@�$�*��$=+����~|�G�]{�K��8_�J��W��k"��i;�r����/�����#�<y�����팖v��j_ )�S�9� I���~,~�����ۣ�]Z��6S�kű������X������~P'��K�W���uK�/�,3�l�B-�Soa��[�������_������`�ڧ��Moƶ�b{�]�C\y-Ps�I��ˇ��|�؉�_�R4�Q�o��ѹT��rI�z���+�"\A�n�p�X1��C��S�w�,+q��<`l� ޤ0{U;�6���Ig���p�v,s�ry�^����?N��lY���=����,��w����P���W�ǘ���+�U�{�?�����W�|�Z��om��\����\�Ϳ�R11|18I������s�f�;M��Ě���=Fo�N���'���c�23����a�WDmV��~h5d�_IA0���@��ek����rυ�>3����sx/K��
�m��#�m�nz�w s�+��x�Q���j:ƫ��!_�)��$�	�k��-�5�D�� �y�W��Z�I�X�aPo�v����־F�G��~��R�.H�;o!VX1�=�Zm[BdjC����:�:�z=���a˻hpx�s��>��h�~�����z�����=�G���$����~�|=�>K_T������h�X�w%K��ڤ�ǅ4O��>LZ���-���ȞYÕ��*��Mm~ĕ��{P��n�a�ˈ$K@�ќ ��7V~�	��o��,�Ʋڈ��r7==q[�_
jZm���ͅ��9{ϵ>^h�)��)8�Vu����u+[��}CPYU��ҕ���F㎄c�\�K�>I�?�aN���c�9�qI4�8}��P��sw<{g֥h�~SyB!�����=:��ʐB�$�!�I g�s�����6�Q�ȸ�1�����-��n��>?x�I�0}ɮݵ?Mao.��\�%ݚ�r����G���=H�k��F�;]X�=��F�5S-�#�9,H��)6쇡������j��olob�(�G�23�_Lx��
㿋n<0<;�]/P��d�����$J���7��̺��7��:h��m�V���.$M�2���=kꟊ_�O�o�/�	���#_��T��O�BrF��r@�`G�ҕTL6:��ڳ◊to�y#�.�so���^��,��,�~�!Nd��^��/ۣ�ŏ�o��t�N�\�K�X\]L���*�/�2nPz��{��;��NM'C��� �5�h���qI�h�ե̩��(�����<x�k��s�G�O�+�[mg�~.��ť��mr�� �(D��e9#����X������(����I+)���k�9c�$pO'�k�,~�2�������������?�MKDЕn'��{����`���B��T�C��*�7��0�ú������A9�ح,����q����� �a���?	͟C�`?��u�?	n�P��t_�DR��㽹��~4h�X�=�
��ݏ���{��� ����7�D>	�P�dh�%y�&��xj6h����G������Od�I�1�����Rk+X֯��N�-m�x���d8޾�q�
�BOWc㚸��&�qm�$�2���W�>�ҭx�x�4V�;���y� ��3Z�Z��X,���1!�Q�îkȼ{���&�4�Oi_ZǸ�K)�+����+��c�`��YX졅��Ҝn{G��-!�Y4n��#>�?n��6�w=��f��ގ� u�N��W��j��� �[O�N����׃��� ��m���ͤ/so*�I`����*y��<6a�ƫѝ�[W�Ecy�&0H*H�J�(�A��:F��^jq�����tm���� �j�ƌ�4v<�^��N�.���O�Z��c����f����;�8��|�wq������&�/�i����G�\�q�GV$��I��m�F�����L�s�D�abl�܊�JyD0�F71�=s�q�_��D��ͣ�|�7«�m/�X���i�A�=3f�&�a��k�P;�%˄��*�
x� ��C�����3h�����Y��9E�g�;�F�9&W�^k�M�Q�,ʇ�Ѓ�M[���<}���ϸ��R=�D}�� E���֗���zu独,㳇X�QV�5U ���p\� <g�1��;]���S�猼D�V�<�o�-�PmU�g8 ����U��3cnH�n2��q�k�o�&=卟�������&k���*������%�RJ1���u�P�=��o,.-��.��`!�E!}k����Ş��b�ym�#1��O��?��^��wZ��rSF�^�4����r��	�Nz�k�'�����i�^}��6��z�:�J�-L}C÷V�O��	$ R���O��wK�.�f�{x�Y'��FX�xǦ3W��V9s��.�U���#��]_��;R�d�%/e�I���B:a�z橦��ʳ�	8+�xN�a�)�G��q ǘJ`:��A���
�&�1��J�nخO�:Տ >@������#�-ꑉ $�èn;נA-��nm&����FVݏPOj�+r���q��|�M/R���^�]�
�6���Cи;c��5*�G$�1�Z׋j��f�}+-��:��o*��2n,�H��}w`�������pɻ�q��}i%��!�o��z�a&�s�/��)Ii��kI����>����G�j�W������.!�+魤c�LW�_�4��ܞ9�&� u�6����E��s��m�9~�QEj{��7JZk c��?ʾ0�����h;}��_g��?ʾ.����\�� ���XV�>o=� vG������9�q�X�"����c�%#h}�m9�?ϭl�J�M�Fr�~��\ιh[E�����<��8�y��%�}���6��6�r�$���r~��W��c$�F=���f����#�9��+��?0��g��DU*���m��eQP,Q�g�jvO�����+y����m�޸��4���1��ӭA.Ia��"����ڢԵ�/7����B�y����n-�)ǝ���/��+p���l��~���K��Xn>�3�ы�b%Hנ<�����n�P��V�kqC�2P��#קz��?k����[W�*=m#<O���r�����9R��~G�P�Q�*��o�?�޽�x�[��!]���kp�ev�d[��#)�=+۞�.kb����#��s����/ڟ�5���5y�q-�%���?�uz.������ź>�ờ</��7�2�wTd�C�ýy���Q��3�.��G��_���9��~U5��z��U%=s���_6�I�KY�[Zm�b�R�U�L���nn��#;�:W�j_��ǽ#V��u	Z���V�x?�a`���x�J�� �1qi�E��&�G�wW�}�%��
��3��5����=O�;~���{;t�����o�S�h}��Aߍ6/�r��2o�9`�yj�c2��:m�5F�)_G�Č@ki \g��_I�I|ls�1 �������o��E�I��422�> v�	\��1>�.M-z[�r�JQI���|#O���[F�#�#��c���s��!�$t��\��M.� K��e����f��e����k���$�`�����_a>jo����'0����d�o���!��J̬Ń����s�Z7�o��4s^ʧ� ��}k�1ا�m�f�?剚qǻqҵT��dpG
��v���o �P0y�(�In.����W7�|Q��bھ�+���|�~�y�+�Z��:��|Cs�*��e�/>��yF� zs�զ��6��7��_��K8!rT�ќ�򩎇r׀'��&��x��Z������I���V�!p~���ֽ��O\_=������5Z=Q�2�x��=)*.ז�O欎��i/le�)�KGx�UA���\��!�4z��7������$��c��֫O���n��_��7��c9�;��J�j�F�㥎�R��	�I8ݷ�/$�u�mD�= �_W��<�íū�wo��l��F�p;Ƚ��Z�O\��CK�;I�N��b��Q��?}G�\i9-�lN�U�u����1[yk�Y]��Q�}k���&��^Mi�	�x@�ő�ӭR־ Z<Zh�1�c��,e6��bh�)�2�Л��{W�� k~�3q�T��6����eޱ�lbrp��𪟴�Ŀj^�{�6�-o��D�� �%#����}�̼���?��N��&W���H����J��O�ڧ�_hv�xJ��K�LuI%W���o����^�0�5u�����N�G�h�a��o��Av�]��b����>���e��M��l�k;>��s��S�^��cg�� ��{ą~�}�M�<�J��)p��O=��`�D�!�I�q����э6�c���ژ)9JWM�j)�)�ZM�r8� 4m
����UA`�]g�`�n���1Z]r�6��0�J�vA�s���P�a*��ά:��=I��$�/���_%�BZ=�w��z;X�G�]�6�3 �	Q���G�7�T���:�C�M�4��]"[�M���;����������������|@���$�i �'i5�g�+����j��"n	�<�z�M7���b�I�fӭ,#&W!H�T? ��:�5&���V6�j��Ѥg��A�nF+;ė�g��qml��1�2)p�H9�:����jZ�O���� �|9��e�Ï`ֿ�S����\���Hq��Fxb�,>�C�z揬��k�-��1��B�Ϋ�G�~�|�}G���dU3�i��Lk���s���$�����۰����Ns��x�\����_�� �X&���A�w�k^S�����͊�{� H������-�xJյ�oY�U��V0]C�H�ዌ��\t�������w�Ǳ�u��n�r�h�� �u-�j��T�@_����^��ψ�^8�����-Ѥ��o� ���^+y�m�ch����	�R=��w������㖻�`(�"J#���S�W�^�_/�>���>,�,�ɯ��5�zB���#!�`�<�|mdL~*��yP���yn�?4m�fF��$pH�~�Y�ߟ
��ZY^k�<��
��\�첰#��_��杚�.������ m��z4�r;K����^/��mݍ�T���޿H�=~��������t]"�Z���k/u��[���gS$� �����[�W�5�u�s����������~b|�4��@�޿�${`W�C�������.��C-������Y��?Y��'�Z���m47z��}��ַ��_Y>��e6��O� �/Z�o��
5�I�i�9��ˤ}�)���5#h�����X����z
�!o��L����{����O�Ğ#F;|M�)#�Y�����W&�����~����u9���V�d��=���
�z���#�`~Ӟ	� �7� ��?�/�^��cDs3��z�l]�f�ӵ~P� �I�%Ax�X+��:RO�,k2He�TOs$�r@���s�sIF�&����9>Q�}܌��;�:�p�y_v���p���ԼM��s����zn���mh�6fV�dԮp27nr@Z�R鿴ŋo������4[���%��ox��I
�Rpq�$p{
�Ԧ񖱤�i�<w�E���j,Ac�
��Hlci�A�g�vz�ý�P1_�[x-tԍm�ĭm>�?�G��$�(#?x��_<	��~ү4�f��SΒ�S�ge'�-�� �=	�3�(��O���#��Z7���j����&)h�ӥה3�n ���?��1��YzEĺ�7�_^���82iL���$���W迁t���h^>�.���)�..�N�C����= ���f��ׯ���'Di�����M�[��kj{$h���g�-e�tǻ7WR��V��ڤ�y'�+7P�����������%��y/�D�I�{����B�������/��OrT�8mw��~i����5��<Z}��ukr"���1�H!��r����%	�����������5�6Ba|��)`>P:v���h�h:�־}�ޠ�:����c`�XG!+��v���/4�M��E�am3�KhCAv���2:��9=i�2�f]6�+����y�V��v���
�^:�Ґ�0I����d�@<���2H噎$#q�t {�#5��դ�e�G�[4��^�:t������HM���BLÀF��[�!X��m?R����{�&�k�U�I���£f�x= �wZ�Y���5��8�QCj�W-�I'9�*����e�Ӟ��)�=���0L���#��T���f��⾸@d�,0�8���3�<t�īG�_*th�$F*P�#E{w�u/x������|!uu%Ɠ��^I������BA9%O^OA�ˣ���D_����t�9<G�<s�����o��`��N�b�̚�	oe��<�����׊u,ڹ0��9��V��A����ƙj�ͥ�7��En����l|�H�]�8�^�g�V�����4�x�>Z$+4׈v��Rprwu��UMF��z��k�  j����n/�#����i�1i(�p�pzt��M~������x�F���6FLGf��d�e#��
}1XJ
ۚ#���G�����;�z��u�Sqpֺ��������<iѶ�ӂܜد4�.6� �M�Y����?�zg��:��o�������vd�J����P $F�݌��^c��a���E]�3��U�Oݱ��g�gŽq��>խ�o�\xji�Xs�[��5��vV�5�mĢ5'��5�_|a
�/��s[J�+��C�pǯ�g��!6��D�d��_�p֭��s��G��4qF]�P���s�^&ͻE��A���c���N��REܯ���>��4�~�u���4%���� �ڿK�Wh��g�q[�Du�c��C���(���x�5���o�����n��H�dhy\���?Z�#Ռ:����K,wr Vs�; ;� �{'�{�mW�p�i"�С�B���y�x�~	�V�#W��3��(ӥ^�_�c��W���#'y��������G�2y<S4� �2��t��T����ERʤ��~9�/��,���ĳ���5�+���m^����5WA�?��&���,��t��%�ΐ!O@;�e�g���4���գ.~Ǯ'���l��{y��7!�4'��5�Y�[�U�6|��ݞ�������]���r�φ+�l涕�6+U�{W��#��{�������m���m^٤V��[y8��D�	=r��w���'�f�� ���h�H��ǈM���Lw�f_���1�����.7�;�����jl�[�1����,�@�[�� ��~-j#���ٺX#��nd,��9�c�_�q$asI�eo
��_� c��|�;�����t)�}]cv+��ۄ�-�s�+��]�/�3��|I��3�W	<_c0�G��YΣ'����b>a�����A�~���h��߆z5�z_��}"m
��m"�G�b?v<+|�'�b�7����O�^��<G�Z��>(�h���<7u���H��#�bTr[
�ȯ��-��Տ5�=�?�W�����_��\jwma��$�]��Gā�s�z�+�2i>����DY�+U��<��_K���IQ�vUI#���k��1|!�!�]|D��ŭS�>��xi�x!����(�I�qe�tG'*O��?��F�D>*���&�����k�ɨ8k���u��:�Q�R�.����O�������Ȍ����Mz�Z�}K嵶� e��w��p<vM�}f;s�Cr�B�)�b���7Z|�6׮eEeun������'�o�>1x����s^�9�&`:�8��R�� �s���������sIXH���iZFU<�;z�^_����'ŏ�薶s\0��y�� �s޽Kş�Rx��=;Y���u��%�?x��r�r�;�.�R;�ٿ�������B{��vx/���g�ՈR�>Q�9�c��
xvk�������,��o�/ְ,� l�Ze�->�z�Kue�i;���=��o���z�qMy��m!�L��-�Ҽ�(��>z����+�gM���I��Պ�#K�+��##�M�,�by��+۹l��̻ �99�+ϗ���¬_��h��e<u��� ��I7�a�iO��</q��k#��6���g�5��8��L����M�2x_�⭩E���?³���{h����E�d�ܚz�ڞ&��9S���6� ����Y�kV.���TnCd��8���;9]"b�yk�z������{������zӬ�ڴ{w\#����������;h4��k�Lq�63�N>_z�f?�k㏁n5�wB�������X���UB3�9�{}�����Ȯ!��|�,#��^�oʏ��<7��՗�w^�$*�~�o�G��[�
� �'�JתZn�m�����a�B.p8��U��_������:��D��I��?ʾ/��c-�1��x�}�'O�� *������dϼ#��Յm)��s� �U�զ+u ��sY�*I�1wmr�[�P̎
�$c�C]w��?'��#iw�^&�W�ƀ�s�08��������G�t��<6ڂ)#�e1��:t?�yTh9%5���x?kI���j�t��i��g��-����71�� =O�]O�s�F���?�@���\��[�+K�r���4�����m�$Ι��!��J�~Y3�g�L�g-'�P�-!���>ÞMq�dx�wq�"�pq�O5���e��-x�����$ν��� 	e�<s�|Q��glqq� x�$��~�����ǟ	<C��O@�6�Vv�Ơ����O�W��.@�Z�NJ\�hz�0�TT�ђk>*����\ҭ��.�V����A��ze��|5}n���E�՛�Թ�W11�;T��<��E�C���m��6�c(o�5�21BK��*��{��_�K>�H��Y�1͈#��T��68�<�<V2�����}>+�ӕG��Y�[��j��m����,1Z�z��H~�0Kz��uPxoĿ~��!iq;�b�[��sr���0r~���7����lm�%�@�G*���l!$��H�v�۴��'W�뗚R�U�� k��y����H�u�^�ePNJ��##�uS~�?k-,zq����+՜l����� �&��߉|}$QMm�iV��۰_�g�T�?��J��j��犵;�f�m+Q����ңG�y��y5�_�>$�E�|����U�A���k�tkH�>\�,�;c�n��8��/�O�Ħiז��\�ז�ʫ gkYz�0��� z�|Fg���>m��gׯM%-Q��ڃyi�;s�~#�Y�m��k�Ӭo/%��N�E��g���<Sx�T�nu,i6�����]������A��J�|A�x�?�z�5�����4M� ��Ae�Ws1�q�Q����r�g���`�g��畹O�&���[��ӯ�8k{�?�?�$��i�ǌ��#ھ�Эu�|-�n<Eq�-�4�����h��̡���Np�ݒ"�������7:-�ƥ�qK�\���ʿ�-f�Lw�SJ�Br�����,�!����{�����\|��BH�=k�񷌓���f�D����H�",� ���[Y�����i:��Ȼ��m�7@�n����]�#GO�Z5���L�%�g��V���\��z}+УE�RG��Rz����/�vi�k6��Z�����TH0z���=��z}懭��JA���KL���K�t鬋�Ж H��X�c��5�������L|�:ͰZF<����V�]s�^4�i��,-$C�r͆��
닺ћ)r��;_~I�]f="}&FO�p�~_( 3�[��J��z�kZ�����)e�N�����k��~�.��(և���
�g�tl�d}3\w�4�ޱu������,�ppA���m7����Y6t�]���ݦ��G� �^Y �ɷE<��O��[=kãPյ��K�^"��.�ש�j��L��~Pq�������+��do�G�\#��~c�yU�K����4�r7� R���ᵅf�����7^k#�ޏ���m[S��ŵ�.�VS,zd�ns��zW�\� �;3�2�rE>���9��_�|����Z��q)�k(�s�]у�Xg��]�ܲ:�����m���j��y4�� �c��L;G�wy�q�A�U�O��v�z��"7�m�r$���|�'��W+��A���[y�i�0�ʤ��^s�y���<e�Xh'X���d��DUC��'B�!$7� ^�T�]��R��ާ9������kU�V�&�>��Z���t��\�݄�H���=����T���zdq�������Y� f��:��բ2-�]���$�u�x'��|#�\��G�� �5�Ѯ@_9B�Tu5�-��#��&��ˡ�5ɻ��gg2	\� g���W�t�>��,���]���YI߽Mg�� ��O��E�g�u?�4���t��2ێ>q��<�y�ܯ�f_��Y<�i0;y���Ё������W�N��G�4�(х��.!k9�uF�vH��A8�>�o�����(=jI������K|G�?-�>~֚L����U?��d]x���i!����8d��Ee>�*9��Z�#i\ӒH�@�c�Ǡ�y"2X���玕�|]�y�Z�A#;^V��"��H1�MBg�sG�ڟ�"�\:du����B#�v���pI��Y��h�+4����~�I֭��.�Z�X];��(8^=��E�H�S=�����~��|Csk��Y5���K(�o�)���������R?��~�sK�N�bHV�D
Nx?1�+�O��O	���5��3���lv;�3�߰5����=[�n�t�iw:M��	�BJ�|���������x�Y3�ڽ�=���?�u�Ԛ8���iC�\FC�T⼫ő��+�n��X	9� z����M"K!�)3�y~|n�O����м/c�n�F���ե��t�Jۂq��ֺؑ��0��2���>��/�����pl�e��%�w�F��}���z���`���Ս�������m�,�I��� ���_��� �b��E՝ż���Hd���Xr� 8�~d�̓�Z�~�a%�<� ��]�9ݙ���$̣��\~�?�4�վ��'���z�#����A�#�_��0��K�vq�~�|mԾ2������+����^�L������BgY���;0W�ׯ�p�������o�-'Q��Q�dS�W�F�e
��H�G�s���l|E�~�� 4}bM�ᧉ$�5���dӅ�Vcw|�Wc�����,-��Y�z���%֭��{��V�o�������~�|T���4O�i�n��;&�R�:,��h=��=�
�������m_�Z��}��ɣIe�J�U�_p݃���RIY������FMcZ�4_��,��{]�%�֎�ؔV}�˖c����z�<#�_�_���ῇ�#�t�,���M�X�)��m$g�k�;�\���k�8�׋.�ui�e�����X<0NM�d]��8!���\�<)��J�H�E��e�֮��T�N[ōZ��m�PĐ��QIJ�w��}m�/�n�Wx����G�Y���N��9>��>%��/�z�߉<��4	o�4�,�Ws�3�OL{����k��B=/H�d�����^TD�m���'�#޸�c�v����	��kĺ��j��X%ź�I#���b劰���5.mŭ�˭�~5�&�����oV��ʭ喙<�>8!]P����� 
_�R�������� �=�=z�����c�����4��泦x_T��Kf��+ ���ő1���.x�O���O�����_�A𮄣�P��O��x��	O���G�)9%������ß�N�j��5����"� N��K/��^f���r�Ӟ�r{��~����v���	��Ğ"{�U�nb�HSˈ�s��9��A��Yl�#U���x��5q�`j�S�O�̺ݏ�u�D���n�5��ݴf�R<`�����3^U��;��#�K��mE�Y|q]�ydy�`�^E|�xl��>��e�dxJ�����4�1K��/gg��@�U|<c
�$��T�l���s]�-���T�K��Y�d��$P�
�ܩ!�#�9�rO{�'Ś_�� O�YhZ������-eq��k��AĹn	@�MV��y"xݢC6�2!'��=�l�J���� �V�G�|2���Ė��������K����=k����O�ڵ�m�Ji�� ��l����c�=�n柇�]8��l���12^A#��a#���9튱�t��s���*f� g�����>\~�����Z�����	d��*�溏�M,/�Xv�zdc5Cĺ.�7�ow!���ѧ��j�X����S�FR��\�tF��$[	'gq2!q��RZ�j�n��I�\M�E�)'~w1�=?º�>�S��፴mX�|Ȯ53�_S��QG�x�T�uk=�,��:4�$��b(�CH��אi7bm?C��J��5��#��
s���V_�/�����n-4�+=�4W|������3���8|Ay�okukoy=�(�h���L��9��'�_S�.u-��PAO�xc��s��U��t7VJc�M�-u��U��MC$|�!?/�YZՕ����evW6�/�-�$S��C���dӒM�΅���y{��%,7��ON��j4�����+<�U ��>�=��UGq�<��֯7��� �2���#�e��0  �ӽt��M���"�/�u%��g�լYt֓�U����������$�u��E� �[�t�B���Iꥰq����?�KO����[���K��5�4j��߻جC�otl���J�D�_��;��l�]T�<Cs%�6��f;1�%^&t'q��$^�7���r-�����-7O���s/�Mª�6�3�[ia�x5G�g��o�
xL��u߄��Տ���upDY�0ЄP���wlw'��c�`~�6�msJ��$X��j��x����J�{G���-�R?8�?~�7�  u)�V�f���%��6?j�7���ۍ��Z��\��7�w9遚�#x��^4�u���5k��Yon$�ҳF��e�s��^0����v�x�vZ-���O*41E��V�b��sӶ+�;˩�������y�M��,~B�j3��*��P@�O����o��� o���^�����A���%�T��1�-�X��^-������I&�t�c_�p���g�c�`[�Rx`T�X�}6�IU\��\��N�W��=ඁ5�R-=�I1G��f�$�A r*�Ik�o�w�jV����-���OE'�=A���c��*����|��+s5������I�4�Yo&��n9s����i�xN�oR�+eiaFXez{�6����Vi����/�_ֱ|W���tMb+��(�I"[Y�r����8�b�}b��{�K��=�8Ӫ�9o���V���K��O�B�����V�_m�u�5�B{�e��ٙP6pr��)��G��"��h�|��f3���e==���[{���9�w�s�n�p���)ΎTUk������)-�^xD]��L��yܽ��A�[��b0Lc���V���=2��'�Y1�v�\��@�+6�9� 8��G�F6����|)�%e��R�#�|��u�>x�'���\{��_X��z���[1�n�O��:W=�������i<O�x+ÒJc���Ks���G dc��A��o��~����D|�k���X䓐�o�
�����~��B��iZ4]�Qpdy@1П�_P�?�L��ן��m�Y�?�F������-�q9�sR�d���(��� �?xo�V%�a�ūE��I����C #������G���=ń�0%�~R[��w��_X� �3�9��o�63�,q\xe�fRN>	��+�����{_�.�l��$�X�к3��z�c>b&��q��~��?�M]A��~7]"��#u�S��?O����jg9)-�<���k��B��s3DٺR� +�FTg��z��v2�aq��q4r2��׮F8=��\σu�b���g�YAq���c�K�W �y�]���`.�凉�3��)C���o(�Ѝ%��˛H�3���(��N9���o&�,:��r��û+�Nr{~UVk�$��a�3pK\�?w���m��^�-��2=��xU������Q͊��BJ��:���^����̎��乎>���_�	�����-�0����9�5����x��e��u���'�A�+��umG��maycw&�_������9��W?,���U>h���S�5Ѝ[H]���5�y�[٬n���n1�cG5�N$Ki��pu��e�~:������.$S��+.���Շ���~5�-�5�v����{֔���K33�>��Utۋ��e6ˈ���H��i� ���t[~X9�ҳ�}R�WPi�x�?�� 
z����/��}I��k��Kg��P��&�X�9	�E(�1E���n�W�e\u�3^�6�Q�KC�jX���z�s�r������Mju5��d�?����ھ?3�t`u�<?�5}�'C�?ʾ6��b�o���4�/k����W>"\�����Ϣ�Iotr�|I�xUյ�B��X��൚+!p�� ���ר�9���_,�i�S�z'�u٤��2��==
���B����7���xG�N��_A������R|�!��9��gX�7�Nբ�Ú�@ğ.P�	9<��:Y�%j���G�F��*�3� �M��| ��`c��s>��&�?�ש�s^���Y�u��@m�c3<��h��X�O�z���3��s ܘ��ч��:������(T��Eft��G$a�W�	�����Yh�}�'�=��*y���eq�M>I��<�F� �o\w�޲�Z&x	'4�ǬY�7�� �J���n�omd�V@���$w�+���<������RG�	��inu�Y�\�A\g�o��,��*�2UӬ,�O�Oko�K�Q�M������Q���h���0���aHl�� B���|�)$f�9U�-�ϲ�Z�ck���5SK����E�Qq��CpƠ��d�H<r�={t�`�����t�?Q����w�~C 
��?0�8��f���J���(xm`��o����u�O����:�9 1׊�m>�#⇆'�4�V��U�����N�P���R�7���������#�p��t#e�ϣ�+x���;�u���6򉠍4���S�$�Лpq��;�O����?�ڞ��K�J�1\�y�S���7�1��̺G��]��7Z牵�`�/X*��`VW;ف�!q�9�l���WP��[���}Au?|>�7���uy�9W|(<��}�qc��e}��c#:ѩ��??�N��ʿ�tč��T�_�5���u�/�cn]>���s�(�����c���ď�����4�?��Ky-Lc�]��s�� t���c[p~�Zd����ਤ��Z��a`�� Vg$��ٯ�e�žJ|�s��e��rr�t>����5�gӴi���]�� �?��b�����jȿ|\p?�ˁ���� �~A�k�?|S�_�V���Ծ)iA�=B�z���l�frp��Z����,�M�^�<A�jg��$�e.!y�
�>^A�#�+��r�U/g'wc�˳
T�8������%�g��Λj�T�+��r=�͵;8�E����J4Z��+}�1�<�\�������V�
~�bT]K�2�����}�os1@����Sӄ�~��6���,�uh��r�Ȥ��@�#\`�9���էV�Y�#�>�a�Q�;���<�mfy�/.�c��k�y&���ׅ�!s�����C�Ř<R�7�n�[����Hӄ�k|�䃁�9��/Ɵ|}�m�o��� �K�u�� ";�c��,�e��[��ៈ�I�i���2Om�X,�c"`�Gݞq�+�(���RMЍ�f���ɡ��\׵��U��H��N��j7�א1� �z��� �Eq���O�u-{��kx�R���G��z��-$�V��?V�~��^�s��O0��V=0��;v�G��^/��YԴ�F�Y��_nۜ� 	S�;W4���O��I��I�$�-t�Vm?Ŀj��,�&�e��X����\��}.��Ow.C�s��� �ֻ�/�ׄ�⛫�5K�� SlQV!��rN[�x��\g�4��=r��$�c�£�Â	�<�]���xu$��t6|B��Y���� ֺ�=��x�-���\��I��9\����ֻ%��Fޭ�n�9�.����U��j
�4h���/j��jxN��J^2�s䌱9�&��}�)<;����˛��*���k#H�]�_i�j����+��bdbpI���j)�RNu6f4��̙S�d��>#�y ��p%f8b����~U��O[�𥎛Ƨ}�BZ;[u��.�g�^Mw|3�������+ue���6, f~�a�1�~�|��_���6QG{����I�ܨ3s�"2Fg'��^����އ�e�<�*5%��߳o�v�]���a���f!¼��$��:{W���� ���_��۷����|Gm��D0����c�~L���U~6����'�ڊj�"X����]��n <�
��׼c����Z��u;�ڦ�+�+D>U�Ns��kЄ!d}�-:K��џ��|Eu%��l��H�:'A���q��׿k�� җM�~$k3٫���$<t� o�8��F=�2I����z�u>�V�Ĉ�+�N1ҴQH�V�F΋�Zj���j8���kٟXe`�HV
[s�|��]6��b�Nӭ��^�Ӽs���{_�Gŗ��f�����Oz�k�O-d#
�q���g��6�\��9�z���%����&��G�'������?�'9Yc�{�'w�`�� Oq�U�x��������MƉs��j֚��g0�&8��<����H�鞧<��]gß��,�F���#Q��̊����evW����є+0G9���Ҫ��t����L�����6�Չ�i�qIosi�����89�]��'�������߃�weꖉ<Vs��nh�$�+��rrO!�K�h�:^Em4p�;��2��8l����y��+6|�WUFL�W�Է�� e�k�Dw�w:���9=ǥ|� �~��5����SB�����=�U���`�
m
H��� ������ԓ�_����kx�,�Z�F}�6��s����p�ؤt�~�ҽZW����o�q>�O�_5��%�ԯ�$������"wd���}*���5u�Z���v�q�n:Od������G=�:��c�d ��[V�vڮ��+����A��,~A�w�[�حz�����׃��	j>"�l��B�ɹ�����FFJF�I�k¾x���>��m�Y�4�o��9(xb2�汮�3�l�%�6cP9'������~��>(~�> �Ě���6mR/����,Dƍ(��K������{�S�;#�>��q|i���Mb���Gu�?K[I���խ�Yb(�0fb�@qҾ����x:����j��o�i��qX �ya�H \�@n������:j� ���_xSC�4xI��k�������C�;ՎЭ��]�>����oY�?	�[wou	3Z��E۾P"Pqߑ�����5�q����O�)��uKO�~Ӵ;�b�P���M��cp�ħ�WvG
�1/�9B:`�_����ӣ�a�ɣ�$�����dpyw�1�<�5Ei�c?)�|�5�� �g��K����A���fx}uI�]?JKH�%�v�M�� �q�/�>�\����7LҾj����[]=����YXC����aҦ�q�R*���lM��o����[Ok�ia6���[�-�,���H8��8�<�/�eo�?�/�����:���7r�F��Yf�8��!ԏ59�v�\w�e��'��ž�����Oi�NZ����V����:��Dp8漯��;�\|1���K}���z��E��%�2��R"�4� ^R�A��.hjKj�g����������P�6������C�����S�k�#���<�0�H�'�q���s3X�S"%����`��у�db���>�UO �iQ�VѮ+hZ��F���R��y�� g9��P�����?��~1�x�M����7^F�a��o�C�J�����F�5QQ����4W�Y�+�eh�/� �!����u)'��Οg�"'`d>�\)H�z�q��?�麧�>�F_ȱKqo7qB�-�� �}��_9����Q�|-�Gĝ"�J��WOe�uhD���\<r*�,9nk������Ӵo������Դ(�-b��e��#���l���o�y��W�o��	~~��2�=��S� ��I�]��zl�2�^���2��%22C��F~����i�<&/�\L��4��p�����׏��e�:���J�����I���sm|����)[c �J�;r�}k�p�o����Fw���c �R	�1�8<U��X���aҿb#N�3�ec�i>)Ҭ����墂��P7n�m��zw>������uh�5�Ro�X?w1�(�wy�A�9''��߶w�|g�I����-��$��k��I�|���vl�Cp7ܧ�/��u�������_�Dk�I��䳟LU�bHr�r��k�JF��|#� ��Υ��"�����8cv�Ϟ�eX��Ƨ�J	�5)�C�Ʀ��锎�9`�t�PR�������΍��ѯ����v�u����_�9�F23!B$i��X|m�6��;Xr�=ɯyu�9���s���v�k���k��7\u8d\n�ÍF��Z:����º^q�6�8ш4�=�����vS���+b��#h�-�*�<�H��J_�:n0�oV���{���M�@���k�R�f��y�-���iȕg�
�
�V-�곹����`w�T8x��Q�M�8̹Y�0��O��R~"��)F��7*�,	��RW0�[��$�TWbH~@P4��^���=_��i��x 1=gϒ��,]X.�,�%vR|������M�NS��S~�L�p��i����@��@&���-����9"��I��)���h�)QN��&fV�uT?��q��VY�w��w�;i��zB��7���ܱ�{OO��/�L�B�i�SqBX�c%��%�	@�^�,zH9�k����%M$W�W�����j�鐻P�k�9���� ,S(q��=��2_=}</���tx��,n2�#�3w{����Z��K�˽ޗ~ѹ���;��h6��E#糭; RYM�����Uc��[ [u�������M3s�?ݑ ��� >3ξ�� nӕ�=��RT�_���?�������]�� �֖	��h����@����������<��H}z}O*L�2�p���)�1F�Be��F��g.�y��o�}<�>�1~s���Sn�c��4u�p/�A��b��AՔ�VL����E��D�"����T�5��$U���KV��&*�uq��df��4��>���SG�Y{��Z,��7���i�?�8�v�IH��2ao��k�W�ARӳ[�v�,��v����3�t@�䄯@��	B�(L�_�Ҟ�[ˁ��j��k�=z3y�B�D|�0����!�z��|D�Ўy�j��Pi���|��}Q}���c��yS9 ���.M�p�� .&n�t�d}�>'oP ߩi�� !ܝ��4!�V�ÍA�b�L�5]���]�����i��96\���9�סw�D{��ϧ>A�*�X���Z0�����X�4�x|�9�������}�"J����O�mQǣs��oe(eO�����l|�ۤ�0(��$��וڷ��ZG/�z�i��n��~r��m���6�r{��m^-���{e��1�4_CyVt���Ǫ�6>���Ud����4�sa���$]����'�@;��Ě+�=.`��w��w�~���[^�����ϕ�E�zJ��8�}�B��7:�����tq�>>���6��)�e����_�BC���MV�;nե�)��-ɞd���e�{'��w��z1ݘ���g���l�0�/������{��J�� o�W��*��������s"YֆE��x�>�I�G-��\"���ta����y��g����/����,�����L����B��m�x_���4"DJ5�:~� ���njT��1x6{���G����Q�D��h�RX��R�_WhȪ�@<eBc 2'��7|���ޘ��f�^ U�dV&-��j�<�5��T��:N��-����fQ�����;g��_��2�5o�S[��'�Up�/u��o����s[i��=�c�E�@T_%Q�7s���vB�2��4+���5��E�Ü�L���	WP�R>�XT�iP5��g����U&%F�3����WD8E�PZ�q���-M���Jy/�j�Y��ir>#�ϣѧs�e<X=�K�k<����Z5r�e;�7Ջ�zN�l�vE�io�rl��P��	MU�t|W�I,�J�
�K�>�LY8�g�8�5!����L���9�o��%�~�Շ���6Kg k��f� ��烫ىV�7�����<���V��N9�-�-�J1�/"�Z��od����%�h��Hˌ��
��(ˏ�Q
�' �؏k�$���=^��"�0>Ж��!��h��h�����c{�}��(_��s�3�T�[�������Bj�Mi��8w�PeG;��S��6���F�a��5e���L0+r�"��8ķL�V���;����FHַ��I�x��q�u� �tf�$6Pz�q���cǷh�c�C��QTv%�Vϴ�!^�´,��XG��������&� ˨�M^o�8�nc��*�J��H����t8jz�]i4�s#����b��J�6aU���x� 'zu��+�L(�+�����.���x�ӊA����jC��>����>I!e�ԶIh��:�,�VF$n�(�S�u�nb3��4����8dq�F@�^_r.����ׯx����S�(����ɗ��3��8j�{W����k���hX���%j�IZ�Z�F�O?i+��`�>g��fEb"?��F/a�#�Sm���go���� ���+�'?�����J����q#�-��������s̝����tΰ�NUB�u�h6e&`�m|�^vv0��Ⓠ��˷�!jm���>~�G��u���@r�G�JL�{�_*��Kc2��- Rg��Z���鍿1�>��9�V��P�[�����/��)w�P!��V���W)�?)N��s'"�K4���E!�X��1�Q#�����S"LC ^}�w�N=Ǫ��FXϸ�X��8y�>VwJ@|��Hq�^�ԍT�7#��j�:����,�#�c�)ɪ��q=:
�Н?s�cC5�n���6�X^;dqU��2�1�-|aBcӑ]��ŹPi�#NsPA�;!�}u��Zٜ|�E�h�?P5M4;���lV��(\V���4�w�_�̋]�]��ќ杩o�ˬjŚ��;.�XԒ�v��
��N8E3S|����#V�@޴wA��+����>+T�<jMX�"�"6���]h�`��(
Yi�3�@f/pF���-z�ߍy��DmqL�Y��N4D&��C�&p���&`x���:&�e�"���/?a#�ǧN]�����~�s)�a�n�Uh�F��JX�-&֑UF��8���c�c$3ܦ���f�թxۆ��l�W#�(�韻9$ђE�����\�cCy���>�	PZԿg��^����zjƞo��Yb�B�h��&Ӯ�Q�)�mkzw�#;=�O����&4?#�҂�-'�^i�W�!1&ͷ �[ n�����lH}[�ޜ��� �x�%
	�Q͡ ��8o@K�:~?���ԆD_+�Y�?�`ڎ>���쳗!tp~�2��60{帮;��8V~�\�O��I�Y�u�N��q�.�,�B�@��y?П��V>���d��W6{�t��ο��&���^�y�z���Wy�>��+�����D���W�xz�Zc`��P��C�Ȅ'�]kȢ���������+u�i�?1���a~�;��,�_m6�#��>N��V�gK
�W���KK˅2���{E�����mR��K�Q���:�Y�[�Po� �o,��`<ID��1��v:lQn��𓟾��~�F�q������j�AuX����͝S�-��>k�W���s��D��q�WV-�Ic@�R�����)�5>����9�=���lY���r�_���4�(��Sx:h����oT��>o��~�L�q��t�Z8�FO^~�4�j�r��6�GcM��Ђ�K��/Ң���ͷ�+չ�LЯ��.��Z0���|/	؝��Ք�o���k
>��yv�2���1�Q���j��1m1�c!f�V�ma��T��b�� ���w�~|�S*�[c�e��5�49�d)�S��.Ɠ粒=?c�Q�C>z&�;1��/�)36Ci����������Ԇ�C�j�gv^Sg#pZ�/S���4�{ę.|��L�Yz#ˏ�t����%0U�d?[4�)�c��!�F�P�S�.Yޞ~��S���ԙ�*w˳Hpy6�K��*H�e�[*ao����}L�g��߾�����D�f��:(�U8wb�"��b#�{o��lۃ�pm�G-�{RXH�/)�N�vV���ĭnߤ@N�;��X_��Ɓ�Cy%�wg��(Y����]c���3)\W![Ig���J�� �pe�tX��c*��#Қ��g�/��x�I�A�p�v�����s�`��n�[eP�� �$z��_�m�U�0��׾��m��r����X�Ȇz\H��Z��_���p����	��f<Y�W���ų�6��#���k��B��S��:�������b�zG�u��EV^�=T�g򇖬�ϱ_���[�:���%lg	���Zu�c_����8zS)��^�h��I�SS��Ԟ��Y@'$���w�:y6o����Z۴e����ϩ�qUJ�ԩ���7�������j��ZS��{����,l��+�?zZd��� ���������Ŵj�}恵��@P+X�`�QJ`j~�\�
���׫�����!���sD1�ZҼ��y��/�J�>KN�ʟFķ�ɦ[��~G�Z*����D?,��H��s���R��;/P���c��a�f�]��\#��P
O��Jft�������/��ܝ��N����Az"\Y�
�D����4���Lit:06n�X{�f9��is���x��M��ӓ���~��y�T�c\@}3R�H./�c���	?�,
%X��=�(�N! l�9*�{���0��T��r��ឬ�:���/A:Ve�ۺ����Z?����|v�\OJmH��u:{Pg�yBq~?����\Q�g�&%dg��_^�c=37�A��w��<�Fn+9������N�W%a/����8ڂs�	h�y�F�E���L�4��`�F��uO�s��{�m|�|�}��z��C�ncW�5���7���[;
/j@I����+������?��;8������b��[l�bY@��p NØ��E��e�	������F�l��ҧJi=ź.��w�@!��- �aMP_���W�OW� pz!�'��^�R�Ƹ͗(��7�����=7cc+��_h������!�i<h��V���v.��D��  = �x��A�GZ��Uʝ�䬦�~��ͧ�Pw4�F+�S {� �H�%S8�o�����̙b�6��\-��u\[��4�˷��j��],j�%�|ӷ����_X���k�FY�N���L�m�����v^� ���� �M�K���Vb�|�Ot��}�LŚn�mC�����0�%�^�9���*����9�����^V!�����Ȏ�G��|x��;'捷ko�C�g!%^�w+"dd���7�-s�6W��1�`9���~���igiVa�""�=��H���
�_�Q��QG^XeV͗v,=�T\{6g"%:�8Q���;�Z��ӏu�%���ж+�3�hg�^k�:�sD=�}���b:���F9����:�@oq�%6=k4Ҡ�V �@�|KJ��MP���u�s��)6ί=�	~3�XNa����GR�S���?�T+�Ef#kT������U��t�0�O�v�fS_�e�h�h��:���j�
2z�Μ�/e�\GO�O�OxB���6�b.h3l�y����B��\��kFm!�'�O��i�/UC�j�I)K~G�W b��]���u���2ĉz��X����,6�2�SE�w3�H,ľ5��k>�z�'י���u��]Y�Y�-O��m��8�-\^��������Uǰ+▌T�
�%A��l	�E��f>�0��
$��5�o��CG����W��L�͐;����i
�:����W[���i+��{����tʯ<��W���~����/(����L	O�>�v�M������5�pY�0?5ZBb�F�d�hn�"7ܶ29~�;4�~����o�Y<�sP��簂����Ă�=�9�p�݂YV����L�l�\��~�
���%��a_�aa��n� Ϙ.�)�$Dk"�ά�F�Xn��;����ܜ�����S/��U/Ϟ�T%(i;�d,u~/�=�3���Ȍ�'��F����-��bv��;���� ��N�ч�}���x^)5@��JƂ,߅�R�J����uJ.��f���f��M����z���2���훂�+����|v�%O�V�:ֻ�͕���������+�W��UE���VY�v\3Ҿ4��4m5�-~Ei�Hx\�lFcɔGN�^�7������E]��&�	�(�w>���4y��"#�����L0��!=".ߵ��ҷ� 7��p��䂩(')��?d���d"���T�vا��z=T�c���_E�@޷%��vaPBDp�?}֣�6Jٚjhg��?�?�M�ȱ5��3 �I4Q5�eBA��^����Dff�<�s#ˋ@�yV22�B����������yXe�6c����{�M.�ʮ��ܱ�bW�	nn꾁K�"W�"��/�=��U�:6sE�n<����}��g��˙��J�&)���+�3<x�X�\���EHԜ3#5Rj�W�be��[��(��5�ʴ0K�B}K<sy��p������'��w.Y�V�e(^1�Z���H=��v��$�4�\�.��G�c�y]�����қږ/������c�%n�i�����Oeg�O�d�v��j�i�A��a�t�G�������*��A�A��c�I��- FtQ2R(�v�#f�Ѫz����&����;|�<�����8?DP�����;�W\���!O>����K���A�ID�G_��W�	_+�8�G��r��,[Ǻ\��J�0?���Z
f>�I��7�$�_���f��4D�L_\K٨��M��n����/ҭ\V��N!��Hl�C���֦�`�&�J)o��w]E90?p(%Z$����Q�z��Q�tЕ|aYs�L�A�gו�_��b�9W�X2Xp���?
.G�?�?�c�a/�=8��<�9)7���N<s���3�֣C�KY��[���`C�@:�.���F@l����y\����,�B��ݹ�>���e�p�|1&��>\��>���-՜��|�i�����`&�8F5�7�Z6Μ��E4����]~�4AJ��a�����_���i8"}*pfe��݆zj�>�į�zrz����r��ePLm"8j�:s�����$�׵w�Gj��ak���@,C~9;�+OFqi	�Xs��#6d����@-]B'�8+�}����;��d�8��<w�Y�ìHA���M{hv�X��L��Co��{9D����'�E,d^�B��n.��hz����L#s�j����� �$�.��X�<��C���������>74%�¶1rp�����O�J:�IiA��,�7�ܙ�\5��X��g9�7��o��A��8H��a�����X�7 �l��n:��ĪqNA4�H�@�1�����-�2^���;�k7#�㝼D��K��"�ED<F�G���ee�T�p]��'������g�6��z�C^,�X(�U7-v�dٖ�|����J4}��y� �%3nPrP�N`����� o��^ލv,��3�Ztz�z�GE|�_�g%��i;�V �W\�l��DVA�ϳu7�M_܌����9�#3^ɴ���q,��-p�r���a�i��������[^�8��q�Ik�꒓�-�`8m�쐪�`��9>��y|���I��fT���s���c�݃��Iv�Y���A���֖Ӥڏ���v��ñ�v����(���߲a� ?"�ޚWb{5�l�l�r�%�Ov��"��V�Ճ$M��z1�M#�Iq�N��7)��	�6�&��4 mE͂ғ��I�����˅�h�d��Q�!e?_o8\8��)���NӬ����loฑɍ�i���.��F_��(7��/	u]�2�\��,��d������"#�)
c�S;�8�D��aV��}��hu	����Ҏ��z��	L:]ⷫ˧��,D,q��(i���_[��� z���LH9Sf��kW�c:1p��I�߾����k�U��Dȳ���7:f���S���ڸb��Le�^�R��~����B�#�̎�H���� �C[��'�j��w�h�Yl�]qM��>0�*����\�j�]��9����k�J ]�G�)�)X{E��E���x��)M�w��:òͣǱB�\�6��yj���g�\XVK��i(�������i���%�ɱ/�j<!T�5B[�;����<����	�w��N\�zE{�nB�Gi�O.�鮺?���%���,�nD��m{%��u�$)2d�_L�Az8�Y=�"S�/I���}l%F�w��(�B�p�X���	������I 8J����0ӝ��!���,��*�
�y�^��7�4�1�	��#�2�&�1����t"1�p�*���S�1@w�4bX�m"���N�4&A4�ie���	+���m4��5�UU�+I�l�6�.�8���xk�s�5��N}O᪚P�ئ�J�oz�n�~��S���7�iF]������!.2�m�NJR6��
���2C�'N�#��vR���66���K�Lѩ0��������-@C_̍Z�{E��;/t�[��J�.���2���㞪ذ��a*��MSm��囅\I~a/���m�<��>�<Ml���uIɵ8F���<��;z���I�I��zG���
"�+I�ON��R��OQ,M�r��7l�+���9�.tn�d�\c��x�h�9�����mS���/�}�^M�W�'�3��e�w���	f���%,�؅����Mw��Ji���7Ђ��sY?w;<lX��eZ��!D\��eӅwP�+�d�u	��Q�l23��f �q(�c<���*�1�����\�콏���n����H�H��t~<;D#Uj��}ր��u�ɣ7#�'؆��?Gl���]�e�bϠU����v�����<˓��$Z�N1;��ο�Phi�����S�K~%�}����h�Ud+d��`�~F�)2����jw�n`GՇy��|�<��[���{����|�&jF����c��V>V�)��tL��L�JX�)��>�Ή�j��/�}-C}����(���x0	�g�m�l�Sv�/CP�N�W~�Ϭ�A�)V��Oz��Ċ͚����ц5��AJz:.V�8�{���'��Ꝏ)�5Q�zF�ʑN��9�nZ!��2��f��9���4�T�����}&�Y�@|��`p|�V�QY�b�20��p��n
��g�t�|�0VVs�J�/ʷ����%L�nG+̬븰�rߐ͋�v\N\�B�Hu���ºrm����ur���3'�^�1���*�A��"�\�W�������Z��:%� ��~3���{	���_�e����hS0O�h�&�?�8��Ū�\2m���	�(������,�\}�A�\�`�����Ju�cicH����?W:��g��E� ��T̀st�gjo*z�%��U�G��.���T�c�U?��y��'N����N�r��I:��M�o���E�Y*�~����'5��Μko۱�&��gx�d���os�9��d��N�ko�|��d��=A�bX�28����b~�Y��Fˠ<��\'�0������g�$(���Tx�Dt�����f�A���[�u) ����A������3��n7���QD��+G'���r�-�|m47hvp�!{E�I�窕��� ͽ'>X�6��R�n����s����L����T�3���S\�l���{r�-����:���Qy�֧��,���5����JCS�7�q��3!�F3���𕽤��M�3��w�>^�& �_��{��꾽k]m��Qw��|W3 h���4�?�veG}Jz�u���˯Z��`�3S=�^�e�S��%�L��c9]�v^%�_Of'���h��	$_T�(���x����ux;ւ���Wv?즏��O?X�+����Lm�T��ؗ6�{��O9^c��0a����Pj�^o�4DY���k�
TٲH=d-5皈��A�$�o0�m������7��:L�@lG��I]ä��?mm[2,A�F��,��:+�p�"t����i�dT��On�0��x[R#��R�ܢb�c)2��6���I���8~ro���4{=��TK��#�?�z� ��|��}D�C|k��SD����3Me2\��-Awu�����+s$f��;.�O������W��~H�����F� '�!�ƪ�b�2^N�C���H�����P��7<i�J+5�H��}��g��r�J�7Ӗ��<�}�s�d�A�����Q�@PlW�c.�=$b:/`6�k�?�OS�(�k]�T9��8���/��=w����<.8�?���~��٬i\���&=����I�FQɎ�6	�%xr�䭓�/a/nR�W���?l"���+�z\�}���s�d�����Ќ��6��_>�{�U��e�������7�A�B��;�o�hiq&� ��f�h���%Z��[_�O6.������Sq�uS4(n��v:���)*q���z	�-��}8v$SI?�t��{�+^p�/�����@��3����k�vM<����5�S���E*i���ǿt��TCV�o�z3�n��F�����0yb샹��u��J�iÙ1!��k`������[�WpR�ԇ���h��l���H��>��9�/�Q)<��߳�oy��xM;�[�JڿΕ�J
��WW�j���U�Wm	Fqd�d.y{���h[W�js.�������~k��s�!�&bW_�����I�����3s��Ҭ,��F��!"� �B��m�'n>=��씅+�!�bvs��Aۖ�3�4���L�Y�h}�ǆG��|
Ȱm�i5�!.IL�ucB1QC�f�l�J�zWӃ!�P�� f�
�p��;��0��aZ�ϒ�쨼��G�tao��u]��v�kC��
���}S:�t�����K�������Ixfӳ~��7��#ۋ����}�;�F��s�ƾ����>�W�O~��P,���{ֹ���z=�V?)A.�2���%��D�ȵ&L���#�n!��S\IlV���.Mߏ�7�I���s#>�?���l��rԻ�9���'� ���.r��o�A��DX�l���$O��À�ѝ����v�	8o'�qd\c�3ÔZ�e��`�������C��;�D���r��;��� �-ʕƝ�i��b�9ڛ{���4�_	�����э��ƘV�]�:q%]�K��Z6S�~��j�ʝ���P�(�s{�bY&�^��&:�R��Xsͨ9���|z�V`x�xBR�H�Y��=.�h�2���2�s@F(?ꂙa��Ũ�o���3q�։����JlѤH�[@H��9��.Yևۚn�(kIt�+�Wfe洓�>] `��\����I粲���ϻ��9���<޷%����0u�`)8��F0{�ȸ1�I*TV+��IP����n~6 ]NNѐY���c�B��Ie=͉cO����@����^A4���8o�r����\+�Nd�\�V+%���EW��n�/�ƒE�k�q�J��^���E���L���������Pw���{l��x�(���9g�ִ)��t�\�	oo���*�+�/���s����Z��t�LV:��g���zH����_u��X�����m����8�dd���Bo Yb�p3���U*��;�v��m�!�9�W�+��pi]�������=�=&hb�J��o�.\)��d'�su���&�7�s�]�����g�`Ѥ-C��+�y���*�<sA���׼��-��}5Ea���ˡ&U|#Ж�p􆵥pya�["��5{cұ�xp�Υ넭g��)��eQ���'�~3�t����l�z�SD�r��ۚ~!i'�����܍j��k��B7�t]������b��!12��x6�W��'p�� `QQ/����ě�r���-T#{X�	��(}�~�7V_Ƚ���rNIp�k^������s9��l�Nv_�d�4׭S��72����v.��S�BH���=�hr�cG	�Hf�sҘ8��W*h�Hu<c��%�C�Au|���v��E���OvZ��ha9G��ɉ��K�N��O����_����MZ/9n�,�=a`Bv�~n�8�L��֞��т�=��^�߶3Mӊs�Q�)7�ZDg�g�Qi���!�~���K��,�^�K �9��ܫ��ص��%����hlǔ�;����93o ���Ud��r����J�\^&���rx.����1Wq�l����5�#�M�LI��W�̇���̟����՚�UP�B�?�T�!�T� [�~¿{�e�}�d)AȂȥߘo��n��{0�F0�QF���������/�u(I�ؠ�vH-'M���W�O�o\��~V5V�h���S`�q��'�LW�"V�|6�P���A<���2a�ɫ�D����)�߭S�f��v
�[��_�b}0;�y "����1��pu�VE����آ��b� G}�DXP�b�즚���nq�?T
�)*+g�t�{�\I���G#��K��8����i��ک�إ���l����C^�"�˞U�#�qh��.�%�q�MU�X���[f��_B^"DRr�=v���(jL�p{ �C�vY_��>>����A���&��n�͔,	�`ۮYq���q�����z��v�3o��q��.�����������.���'������:�R�
���y����k�Y"�$��nә��r�\�a�#P�;��YwG�m��%ek�#ef�9�P�*��	$D3W���Rm
����q��W?���5;i�
s~LW��9�[���,�[�>��=k�ԕg�MI*�'�Z�qM��d�vS��N�_�C�QVEp�0����-�KRs���4�-�]��br>������}�NS���~abCm_��M�57�Wm�� �)װ8i�7�9z�A�S��
�+Մ�H>�������<v�3E�(V_�Ud8U��w�I�0����N��G���1<T�3x�!s�N����s�9f��F\g������V^���5��M�t�E��ngbj���wf��W���8H�=�!����B�e�嬻�iD;�
��Q� С�I�j �L�R�zV=	z[l=bb��x�vϫ���C�`7bf�v/��"����+D6x�Qv3l_}�cwX��q��5ֳ�	5�S�K�|#�SY'r�pQbbë�����1/���V*��<�ga.�M�J;*!m���T~l����'�e*�!����wgb�DQM���Tj�����h��%�Q��)�@��ts����T����wm���:�������R��<�L*5�����hǹ����z��UT6g�0��"ذX�R���ɮŦ>��c����}�!�C�&��}�i�	�������N1G/YeN�Wq��L�7�C��L��)t���]�OS�����,)�G�۝�7���k�)8`&����>k�i�	�l?�ĕ��bEB޴}��\��`�f؋م�n���̓�t6�#Ї~�(�_탱/^a�!]7As�/�K�o8���G<f)^5-|Sc*���O� �QK���?8.���[:��N"�$??��d|r��C���*�G�_��v�~�V��?VH�貯&';:���җ�v���;Oō��f'ϸ"�I��73�z�ID��â�&�l%�"kW%����ea�}��q�B��׍d�Fk�y���2���O�ets��kF����I��~y|#�B��\��׹�O�Rh�|V��>r���}Xi�@�1�,q��g�%� E�9^q��*�LzG,�&D�Ǡ`NgW�5K�'��F%��t��u�C��ŵ��v��D��%�-�Ƽ~Ũ��,��D�R���zq�Wޱ���� j<��4���TFyLo�5f_����_b������>e�8����u��)��{�G}:U�����hiA�i�KQ©L������ �Vz��!,u#���_#�L{g��{?�C�(���Np����)�R��kaaO���t\i[=�o ��dv�ٍ��iS�.mE�\�܀�=�|=�e����%��H���(�tp	\�6��{��1�q���M���vh�X^J�ܭ�tQ�F�ĸ�����_>\l�飊r�Jƿ9�9��z���e L����kܼ6�X��k�)��O�7E�{/��d���߿�N`�`t�+��3X�{'_��2�4;D�T�rn~����Z)+��%�vd("�$=�WإH\=� K�͡2~���Oa%����`�H�!�V�ֈ׍@P.�2���<ݰM�T��<���)r�@���(��Ŝ�K"8��~ɦ�0�[��X}]~n`�����K�}OgZ^_qQ����ޖ�K��"z�9����L��=3�>�\��^iV�B���Չ����ds)�����s�;��n�/�O|U���)_ ��=����e���k���X�$5�
c��e���$��5a^.%Jz�3��p��<<CICm���ov��F�)˶�m�+\���]��ZA*�{�tÂy��j�1)��r)I��f���DLL�`��(f��I�8I��ت����`�/��Y�4�ד��C%�S?!$�B���;3�(��|�U�}ov��WWBwPH��j��m�Ps�1�EL���[���?�e4���⹔��ϱ�KY��U�������|��]U�u��e�.:TK�V�3��6�\>�l��)�����[>N3�����n�V>�G�P�n�`�qͿ)<ç�r��T(TM��5���y`m�г��T�kg�D�PE,T�b���_H������Ƶ��\i1�?�H_��/JtQ�acs /$w�J*����<b�|TS#E@���^� W�LI�����Aú��l6�>_W�a5=ev�R�4��y�G$�+������p8��Ϳ{5��*��/>��۟�B]��D�n�B(�K�D�t�F�nɢ����O&r�ۆ��d���N_�(��!H�yK&���y�"���:�:�dQ�`9߳p���۠����(�:o��i��ٶp�;�81�)�[��q.���=k��5����;�ܘ�+��H���<e\��_$��'����z�y븾�G��p�!A���h�C~t����t�2�N^����G��df���l��I�x$�3�d���B՚J[3���n�0�w�#���hS\B�p;��aN5|�"险hT{2���hf��r����ԭ�) �KjO��XA�cn�!a��(���1_~�O��0U�������./vX$�#	�x���mGo���"�k�������S��;}Hp���{��qGS5���c*��-�mZ���� ��Y
�5���[ ̙X�P�#��?�����ʻ �u�xwn
H�r�λ�7��Fbr?���橭p�r�b�KnQ����XBD��X@7��/"�����ٶ�8ݍ9z��W������7�b���^>�� Q�x�6�-0���C�K����MV�'߶=�c��n:|)�:���L��h�6c=��}�fu�m����T��~������,���[���6s��FA��\.�u��L��Y�$���+�S���&B��ϸ�����պ�ch.}��R\M睬�S:�����s�0�`�����Pfn��H��Q�͈t�q�&�݄e��d�v�������TY;M�%/5cn��L�-�� F��E���D=n"��Lг9�ʉ�7vW�9��9��
�zZ����ޮc�JY~x�S��Γr��-`_�;�:����
��\�d�!⢸����X�>B��>$�(��
��M����σ�'1����1���s�ꪫ���8�2=�A֣�hr`� ��b�ޥ&���jH��=��^�.����`�8��!!��F���s�կU��b��,�B�\�~���k��uv�K;fC�����wq�U&�"	_��u�.-6�%��L���%ԑ 咝߯��X,�^��7j½�u�i'[歞�;� F<u4eC�I�uWs:�ĕ��q����ͽ�m�D���H��+�Y��R^uI�����s�bH�G�ZseX�+\oߛo�+���6-1�O1 ����1p�Q6Эi~�;�O��)O84��XS�Z�]^Y\)gq@����)נ��<?��oG{gkl[73��.�����q��ֈeښ��ѽc�c���c�Ֆ�0A��u���lJ$#���+�h�J6�3I������\�F9_H�Ra�ӃX\Rh�	Z����zj��Pi�}�ˀ�|~P�����j_��΂�Że�Z�(�)r!�+N�<�6���=��RV���d@����Z3�N��'׵5���(?y������|� p���\q��<9C�5'��xST���$x?� i�ece|Fַ��6�=8�Zn��j_	uٴ=n}=���pzI���S�<M,��i∓y+������_^��������j�[�la� c��IG�-ߠI)<u�[{����i��%��7��⨼<���p�i���=�`oت
�{�sǮk�ࣾ$�ռu�m
�Da��]A��s3� s���}+�� d��R�_	�A�j�����`m�Pv)1�V^~d<����� k��Z[�Gv�M�vr�n_0���7W~5`�>��f[Kc���ai!�X�N����-�o��o�Y�>`P���?3�u��b<rT{���C�{���;Z�<�iwb�8��7�v�rv��T�:Ƹ����?Ʃ|3ة�88-Y�f�7*I�jv�t+���r3��Ҝͱ����{� ��fR��1�s��}�C '?1��iWu�h�e�w�����Rۆ>Q���,o�\��8��eᑡc��鸞Z���_]�CbZ����d!y8R_�c�9�H�Y$��P�� �_.ה�s�O��W�����2�~[�cM��*�g�L���y�(� �ƂQ�očI���%��׹b�i�=�6ޛep~����՚�~`�G"������� ��t,�y��V7���[<������ۀ0�h��M1�|�T�4�~P��Ӧb�;�*��`�zV�a����NV3�i@�)��Pc�}h���z❄n�?J` �ڝ U�84 Ы� �4d2�G~��#�}qA�� �'h�ƘPy���YO^���''ҏ�� t�y��i� uy^hPU����2qҀ[�WԘ}�FQ��jזv�<g�U�S�gK9*2W��NJcG����|1��'���W�+� !�V�� Fr�&�_���l�.���f��[�q{�h��e���m%�8��#F�N����C���� �� ��m/�4� Gop�i��̊��8(��+��?�3�}� �~��m3��0k~�y���H��������7fڽA�q��z�E5�����Wÿ�Z|�i�+Я��MMu�8�`�dr����<�GN����ߊt�J��/�'��y����{�uE2�K����*�I9�	���-�����	�hګ��� �X�u��G�#f�d`�q��rqھ��w� ��M���/w�����WV:���k��u��<�{P׽tJn��>`� ��j�u��O���ՂL!�g������q���8��T� �x��!��6��m}�K`��>M�e��+�m�<w�s_�W��⧀4�";[�y���X�FpzP������	����3��<k�(��3Nן�PޤW��D�H����e���:}�[,|C��|����a�
�O[8���5�+l��0��@r��$z��ڷ�o$:�ڭ�]KP���%�B�b4�������$���"�G���b�⑱�^�#x��"����rY˕�J��n�py"�.�_�R|A����mWU��O��Z�������!yрX'��VT�{�Sݵ���%�,�:��me�36�7��;�
�����%�)���v�����f��?�O��}�ۭ�����.��<N��!R�7��9ϵ{��~��E���|Uৰ��.-�x��YhL<�_,�Q��:׍���Ծ��$�ǉ�Ye�k���2�qoz�<��D�F��=��a1�wf��j����Ǎ �-�4�"��Aӷ�>���|��0� _|��� ��ů��c�]����UH�?͑��1�ǧ����$�Fe㜀z���Aȯӯ�%}���?g�>��-����U��<Ǉ1��FL�Sp#�~��vW1��8�~���~2x���M>�A��:=���0 V�黷,}+Ȯb�����u�=��r��T�&0�I
�6 �A���{�6�⋏�2�^/�K��O{;�I�}���l�>f���~^x������|A��Z������;P��YR����o1���6 � Vq��\������	��{��Ė~��5��/C"_�y��y$2�A��&x��ǿ�J�kڈe���n�n��T��UX�� W������w�����SM=�9ﭷ΄<�#�n�x�+����o��w|9�Xk^+��;(V�+au3�+��G\3���N�$��?,�-�-�3�4lʸ�ֻ;�?|?�_i�h������?�BvH�3��(��'�Vy`��7q{,hex��&`��}��tq���暫� $WO��&���������D;9� 
�'�_��,���HG�B�G�y|�i����i�#�dH|�U-3a'�6 Z������xW�]���]G�ƾ֌���k�6�T�@6��9���/ٿ�w��|U��>��ø�y���� �['�ڻ-7�� ��� ��i�e��(�[�����(�#W�r1���9�jȸ�E��?¾����LM�5��m�N�Ds�9���I����q�������}g���c�_��Gh��;����r �}_���?�'³se�X��<�������Oi0*
��|�A$�o~���|L��>#|{��N�fѧI���i���2x�I�>o��^��)��ί6����o�|m��w���cػ��D�|��>A��f��ڣþ1���gӥ[[��e��6���/`�Knt��ͤ�n��^KΈ_�����x�J������;�//#�"���Y�yyl��I�m�/�O�'�[��R�|?��֩�( ��]�� nϹ�gԥ��mc'�o�/��]�S×~�+�{�˔�@�� �%�8�k�#�G�|P�?��C�Z��;Kt���XI�&RKs�����m��|O�Mz�K�J�ӼD�)���Ir�.ݧ��G'>��������S�4oiZ��/�]��~�u ?}�j��F@�2N��&�EOM�� �
����~��L[�=
��V�Gn/!��iJ�?xdg�|a,�Lb@�sq!	�]�� �>�Ҿ��?���G�b�Ń������	t"��oI摅�8�o�>���S���(x�A�� 8~A�=�9��T�ʵ����'E��|>�;��ng�u�	<5�d�1Βm�Sm^O �T�+���������j�w����s\i��G�f�ޠ�1��m�x�H�C��<TuVK�F�i����r�U���,O|d��9�5�v� N����0^Z�mu����;�^"��Ͱ�}ݹ'�ne~�;=CB���a���\�����[��̓��wU^�<��Fާ5��$�����BYݘ��r}�I]�Y��F��o0�#f'������q��sH��6qQ�s)���;��+��F}h+��րct�/Jy'[���08�Hc*H>�*{�x櫽�F�W%U@�9�[p �2��>����ZD�.-��I��r9�_B�&�%���_�[h��9������p	 �ƽ��~m�MMq��D1���{��ϛ������'�VVP�5��H��zV���v�VK��- �@-��1�rA5�Z���b��/��F����M�kɨ�yl�αt�dh˨ �ʉ(�qjTj�� y�,åR��U]ï\S�V�r	�x���T����;yB��%wc��ޮ1_�@��D�7^?�U�o1��`��ˆ��#�}*錮�~��l�qӿ�R�J�3�o�+�H������ �qW�_3~�<�����?��U����z?
?r�� �i���)��QE W�?�������C�Gm�M���1#!"d�G ����x���\�l�I��`����e&E��A^��2WFUi�X��M/H��%�iv:��V5��q�����3��zū��PxZ2��nKO���T����kIռ��Ig���x��௓�
�\�u�5֛Z���j�6�_5�)��{���/us\�<p��wl��d_/`�9Q��9��"�(�\9�,`�Ϡ�'�W�K�"�R#��� 9��f� ��7�O���{ۍ�T�z��N���f٢�(�I-^ǃ��3�1�]����ß�n��xcR�|Ɨ���� �+K����}�k�-�iivS�G�-ʑ��7��,�I%����(� �h��89�~��q��W���~�o$h�QSjy�s���ھC-ϥ���*C��e�p��P����c����f랇��W�4ѭi�6Y��q�p ����4����;�����H�m�Pv�7���y&���?*���f�#�׍>���V6���I&� .�1Cg�^A���D��|J��Q��f�%�2�F���+s�7���$x��K�R��;{s;MqH���u��π�
��7�� Y�0U��j�c�����:q\�2�2.�"�׮��e�������M68� �� 5��-����p�n��<ƕ7g*������^������>�wW�u�,@�Q+�'�5�߲߅���Ⅱ����|������I��5c��t� xu�t��|vM#�yj��p�v������th����K0�Zu1���%�~�� 5-�4�2�+y	e�8�,*���)|^�KDm���kF�����$���󀻰C�W���}Ep� ��+�;o8���b����/,~�o�EXۣ{���O�w#��z��;{&��sȧ��I[N�m�O�������S�V�/���%F2F<�'�}k�/	|v��t۔�f}�D�j��N0A#���>����ڇ�	&�G��~s88�̞Ƹv��tMĲ��Ð\�㷚�0�@s�\�������gn��%����V������؟��B�Zpe���?�U_��\�ȑi�[��~��i�ֽcſ�� ��+���^h���m�K�=)$C�%X���G5��ü��6s�+���p�梏?��xi8T���c|?�������Z�b����.��o��RO_�w_�7�]gX��&���w���On"kX��d!�a���Mx�ŭ�&�_?9��W��P�w���g���zG����!H��Z�P���׿JP��)$������ڽ·�g�;o�_<f�O�R;� 
��Ȗ���Kq*&�#
s�N	��/����^�կ�!{s�7K�ͩC�$W	�E��p~��_3�z����Yu]3S���ԓ��.f$�r����޷�a�s�=���^�=��fJfդ�}� ��5�]5���Zq~�-_C}"�5_�}d]�3#�[�>�?]�*�����ֺ�E#[ɭ�r�]ftn���~/����o�9�(�|���s�l�:wɮ��;'�cHf�E��$�ren4���R��GN+�R�Sj��Hb?x���>��p�͈�o������fO��|u���{����i���� }�P��S����H������mv��aw4ct���8�O=}����'����zm����o~Ռd��ITө�?��MCC�U���U�tY-煤O36���?�|���F���K��V�.��M���|�F@�iQ^���J
��i��	��:u�S(ڡ��zrWM� �6��4�6_e��_��ZX�G���e��z��4�#�r*�ҍ���-�h���Cr9^*V�o0;6蛩Q��V�5e��I���O�J�dG�"�hY���ǜ��l��Z���"݇?���hAW'z � �}n�[�YY�:�Ǧ})�7f�$QD�.xt޼���j��V�}�ު�z����7:��8����A�c�9�#9�ۭ6k#a@���4,���#���i�pn��jښ�&4A@'!U��,6j�����ކ�q�F��LtS�ը��U+��g ,����W�K�I�\4L���q[V:zC1m2�k�Rs�P��Y�h���*z��� =k��A����9n���u���>_&b�$��2�|�i�7��I�6�3gs㎟�I�A�O��f� �T�-����A�oA+�Z���mX�y@<�W�_/,�� �\�<�[��k-�d��$l��`?¾-���O�7��� �{c>��SM=�	A���L��? j?�Dqa����A�<�jkj�UR�.GLq�q[�̙^{�����n���z �#���<����|�x'i�2G�ϧ�Hl�r�Ф�Ob������vیg�� �RJ��>j�{������+��D�ˊUR�rz�n�� �lg���O�*H�lĤ�%���������'Pv��z{FI|�0*� ��8�� �c9��2y��afr���@ {u�=)*��������,\xż��2J
2��v?�hi�$|21���*v`H��xn�����C���1�!1�����@�� Jr�B�]��'��u��O��-M='�Z��ui%��y6�+o���	 ddz�W�k��5xFKM���[7"�Iy���P�.��v�C���\�x��by���t�(k�	�]������~�c(�9�a�����)XA�t�綖�;���~�Z_���z���$��q�g���A�#9���mM�_F�O�Mv�"@��f`rI���׹j��5���u;�;�k땺���N��{�+4YU����~��߬i�CF����q��# r~l����+)=Jrily�Vg�F�w��$ś*9$~�����L��T���	��~_^�����Ӛ��d.c�T���>����̧�3���)�_�����F-�'��d�B���l#h�x���b����9����Q&�9R��s�G�<c��9��Hb�
�?x��{c��G\q�q�׳?�+5֓�����v�ב��Np6��/��� �ol�-�Q�x�r�ax�;��U������
9#t�y5�>q�b��^XC����s�\��,�9�O2��w8��q�J���_�� �|e��LOɧ�lV��^7��v��C!��g�� �H>����-?TA[�bRT|��p�G5�.��7�?>�P�{PM��y!���$��a�XY�\Z3�[]Ìe�q_��� ���-��!�����k��.#�[c��	 �����k��#ཎ��?��b;���Kb�������q��{��%�R����%��I��(����`ls���*3
��[u�m�r0/��h{�ӟ\��+�� ��|�P�x��HF�D�}�x��
)(X��q��'=+���� (�G�#�6Zn���X�����-��Ȫ��[��H�ބ��n-�����$��y!K&�x �p>��P*�L�'�|��Y\�낟1�'���%�/�)��xn�I��ֵ�a�<����$�
G'��:c�G��'���o�|I4�������NF�spћv��.@f+����F��|�����#{��ˉ ��Y����s�S�I�h7�.���s��̭!#�^p��)�s��`� �j>�t� i�W!�I��<���݀��=I��k������֖V���7l���}D�
m�*�E�NA|��ܝ�;%u�󄚦�ۚk��\e��� w �)��0ɹ8�'��&��Q�����Un��<o2M�[��d���϶�ǽ2O�p�����%�1�����U��7�On��(��#��'����<I�V|9ӵ��tۍCku!*X#l��?O_���_|_�GX�Ss�KMcY:{Ey�'�%<���/�(����:�����v��?i:텎�p�]к��M:�6g���d�0w=��� o_�?5_�V�>�=�������C�۰"L� ��㞵�\�]Q~�_<e�<��	���מ[}i�D:k������&*1�㑑�A�o�
	>6���2.���_�[�uf�奉�}7�g�}+�<;� F�=��Վ��}�r^Iso�;>�K( � ry�q��omg�w�4����ԚT�&�ł��U*J#��2A9�~��Q���}���x{↏��Oi}�_fOIjN��~6�
�<�W��:�$�S�T|,T6>��_�����R�{I&*�ɒx�+�/~�W����7�cxSAK�1ͨweO�q��A<O^k����tD�:��B�}v�k��-�1,� (���\.�2 �����W�	�����c����KRд�&���0Y�$3@O��k�� ���>6~�~4����x�S�[>���t`��@�nv�H#$0#�1_ |��m�^��m?�Zl�x��H��HVس6��P�6���ڢ�C�k���~(𥟂4�KN�V5��S{�T�E��c�8Z�b��� �.|S���w��f��� �]?Ot�С�m����>�%�?2�䜨  k�����m�����>��{��ֵ6]6�2�	Q�܍�rq�N9?ak_�T�x�B�еo��~��[���˕��YQ�h��q�z�{��o��a�h�-�MSR�k�3R������ QT����.�c�6��Q��4˫K[��.���*\C�@�Klu,�3)e`A�9�x|�qyw%��Os=�$����S՘�:��)g��T����W�i��nf$��IbI�'��������h�vF[��<�9# �w t�r��y秩?��rI�#�R���Hm�ǃ׎N~�)RTh�g�O��E=����H 
N�i��u`�x�������b3�q�<��ЏOqE�#���兛��9�1d��Fṛ���y�*i"���6�ן֐����F�e8Ͻ{���UԌ�C4dׄ����n.�k���� ��Q(A�y�� �3��)Ŝ��߉L��b�W��P�o3�R���5���X����?�����:�h�����y�_��ͱR�*�g?y�����Dh5 ���sJs�Ⱦ��������,b��y?J����J�Cl�C!����^?�=@�ه��(�e�x�j*�����f�G�R5�{;�t~��?'� ����.*�m{�k��)B���	L��}0����GH��\��ʟ��QEQ�R@^K�FIj���K�-����_/�����Ez�|��nkQ�bYMm�7�����I+���j%���jѡyG�?��5��g�hQ��J�����r�X���ןOZ�MI�=Z�t{�d�,�H����b�g�Xh1[}�/���
4�#"09�9�֯�@����W���v���H����mP2'�ֱ��q��<�OM*OU��;R��/���x� 
�W�լ|y����Otm�;pV8���c����8�J��K�?0`�}1�¶��:��k��:���O8�Lc�&>�<�J���ʏ+�����|�yn#ڽ{�T�;�o�]�%���pM�,��2��Py������E���O�'Gu����4���1;U[��'���<����{T�k3�_�6�����&��w���9���~"�i��9��v a�f�O־g-�ja�0�����>�1�jX�j�5��~ ����K��_\MS]ԭ�Qwkp#Kw`ʸ;�OL�o���&��8������}8][�hr�Ce؎ �ך~�:�e�WR��Is�� j�hWz̭�'��ҺO��Լ	�4�X(�m.IJ����J���3���|#�����'��w�<R�2ƚl���%D�ǧ�J�?c{{M�92¦Ut���˶~��~�w��|M�K	�F=ӷN���~�dI��/��*�c�����g���d�ϭ��޴#���nQ�Ű��+�/�b�%��|�1ˌd�y�U��]<���e@�0:u�|��k0�W��������C',d5g�<E���]>��4�l̏!�ʾ��.m/!�n��H��v6,��3� <P~��j�.$��-�#�*����T۽t�-�r�ή2�ލ��b�������� 8�ȮG�F���+�9+���K=k��f��A�&�{t�?��w�*��nl%q� d��XiK�1�����Uiބ��QGoJ߲6��n/� ������O={WĚ{m�2	��~�J���4� �G�P6���� �5��t��j��&��O�W��%>��+��]�N	>���J^ҟ���B�u[�1=����cg���Ȋ%bK�����_���c��1?��5���f|/}�c?��#���X�P�b9�q���?{�^i����o%��7��p ��w�k��2�9^=j%FV��xհ��o#�!尫��5���GQ�L�}��P�̸�}���y��j�O_�ͥ�<�D	fgD��n#'�dկ�V� `ԴMSP}
��ԕ
���Nm�˹�Q���ܱ����.|76����r�f4��M\0��(��]Q�A<S����B����6�I�����w�e�돧Bm�,�I4��?�C��v�=�ݭ��=��,s��sg�i#l�n���`}zW�V�[��ӋN��ԭ��\��j��g�㚯��.�]84����.����i6��oNÚ�i-wMvD֑�=�ng���xێx�j���ͣ�wugh���~��Fۢ���[�:�k��W;�>����+�j/��3O�(�!��Q��;���jZ�W�'_�$p�%�J�k{�� �8��W��}���Y��O�J���R����F8�����i����K��km[�:�Koqd-�U���92���B+���ғ=���\_�ύ�7~�N����+�<��߮+�4}q��'��f�� m��3|��=�
|/�7�l�ڪ�;	��x�����t�:��=��gut~�)$��ߤ�J2<�Uy)�T�*uv�Y�0����o�<��y����)�>տk�h�*�6�Ɲ�GA4lL`(��=j8�;�2��z�W�(Tٜ�xc�{�M%�Ŕ��+m9�� �ޒFe��S�,�	
:r{гĨc\	3��?^����pě7�}��u��(m��}+L�L��%X|�0�Ny�Q�9ԑ��`��/�H�ۤp�U$���/b�gr[w�尤w8��`:x�;X�"�W?3mw ����+ʹ���x��N��W��UT�������k�&�t�8��p�!����}s�ھ��_���ºT��F�_���|<ڄ�*i�ifE`"�ʀrK/-S)$�Z�����#6xcE�3�}[M�R��nd�C$�#�BU�E8�0B�g�Ep�$����g�Fվ�~�LQA�Y[G�ڧ�e� ��n��X J���v����̩xnmf�vY��F�n�8��k���[=b������;�]Q��tȿ��� ��q^O�te̙�O:��[��A��|/𱵴��&�9�Z�aZ��^r�&A�>���9�h�.�]��~�)~h�ܭ��S�n8>KHwG��ʞ1����,HO>�M��iO�|�g׺�ݪ[�n%��"�c�����ӣ��z>?�g�ʍ�cE��}OV����;��=�����/�d#\c!l��0�{��?>[�V�O��;�]@n�K{y4t�(W�ar̀�~l�� �_b�g���7�؁���?� ��� 
�5�9nA�E�ۋ�M�1�'��� {��KV�pͫ�����J�E��� ��쬳�J�L"6�ځ��r �U5O|7�ƭ���?�~�P۞��#�c`����N̤^B����њ�[fߞ����N9_Jt�.��j��UM[\���KcN>����4㉫%�һ���"��o������#��L��>M�LcR����#�����3���#��S��_�������� H߁�����1Ӿ99����L��Tj��q���T���t�Kh~�[TlG^e��7;լEh��k,ζ�;?��ᆡ����%���yrI<)��61d�|��GaM���>��1��?��Ec���4�[�HݎU��ܼ䟥p0Z������l��WV��?2��1֡��6��f���G�^�L���[s�*���Q��1�xm���`�h��V�T�m�)8ٽ�e c�3Ҟ�_��ZG}�V�T�i�&��/�Wk�������q�y;�&���,�H�.�����r1��گ�i�R��ϫ:���"?s���Cv=x�W���R��u��_�����|:��ݪ��z5w��$p 0~_n��V�A������?��V��8mZ�է�e�����k�Ԥ��N�"���� �ql�.�. '����h:�ޭoe�7��QK�$O#L���]�𧎸����[[�ژ���_xw��oog��UӮ-�ׄ��r~���q��^i�����M��2��(���R�����}�F=1���{aa��Y��g�ͭ�x2���2�y�pFW���y߉5��jKq|6m��5
�FN�8��ִ�V���h�J�{ǣx?¿>"|Y�4_x.8�R���k:�����<�]�sЎ�t�w���֓?¶}J�϶{y��Qo.N�\# A 鑏�w�\h�<�u;��=��K��KN�{�5�ߵeŦ��o|J�?���E��c
��]��6W���wӫ)Ių���]�s�}7��� �W`���!�.� rx� v���� �sl�� �_k��Th�Ԧ��n'���V>�}�y��r��V柦Aqo4�k�!��y�km�=����L�[|��o%7�$wȤ��;U�9�o�[=B��*�h^k��;H�7|�z՝K@�H����	�޾�9�f����Pʁ�G^:t�1���� �If���\��ߖJ���">8��=�ךև�� �-m�<�� ����k���Y����9�f�YK��m�<m)�t ���Fi����}�����G�Ⓧ����?�}:�������hLkouq3,��T��.;�^9���>i���N��m���V�Y
����q�\��񟘬��8�}��;I4��72�`{t���ٌ���(#�m��SN%V���Dϝ�`�W��� ��ޡŧ�+=�P���yN���'�A��Y1�sB�a+Ы(9��4z*'����>c�FA��o�&��T� �7&��|2��V�vOn�F�ۿx���� �ar;�\���7�*4�t�c[�����Q�����#'��Z��v���p2x�R[�&8݁�7\�C;��R���/�6���/�[�VU����iK� S(�<c��9��V��
k{K�3��ޏ�@���<7J9`������$�x��-7h��ߩ(�q���~�z� �����d3��[h��_X�
׼@/�����֒ �G����7��gr�g�s��+ݼW�	�=��"<S|d�4��I�:���YḞ�y$n�?�#�S�G�5�ƾ)�m3�PʷV�b7��9'R�'�^� �x|y��k���5����Nn'f�9Gِ0$�T��gs֟���J�g��S�G�M�xv_��Vҿ�ǈ"�g�x��A8�Ph���x>���yz;�����E%r�3*<�]Ï�����A�'�ۯ�K���X�����čo��� 'ʈ�v[���M�M�����>k�w��=�XƑ��+o�Pr=A��{�sF����h?����wH�����;���s$�*�m��
���y�� �>B�0ZZ�k�w� HMQ��d��9ۥz���_�\��o| Ե��pݺ)L6F�8�<q^;�?|J�������F���}�M�N�e�P�X��O8���T���r�^�3I�o���"�]%ϒ#�V�@�w�;g54z�����EĖ�F��_]2و;[gPFG>����n�y����f�� *�������O����1����������O���io70��j�0�$��T\�w"}�#vϟa����Y�X����Tqa���x��<�J�4/�_�qy�âhZ���J��=@�"F�7#��3�8 f���=⯁�U��[O�I�q�\L5-6�̀T���
�:����^:֣�췶sY^�-�YJ�E�$`6�9�ϵs���LFcV�Mj�u�?c/i�?��ş�����V7Z��bE?��`���8;��~þ��:�7z��Z�P���j?�;�Dʥ~nT���|�]��Z�o�{�~������<���6�z��'��w��}��8�MB�/���k4�}�ᐩ�`0�N(�yӏs�~��x��Y�m�߄�>)��|Cᵷ�T��+ݷ��9Q�'O�'�~�����{��>��^��~3��5���)T$�0Ã�A�?�2x�mPI�=[T�� S&�4���c������#�����K�+<vGV�ً����!���+ZU}�����u9Z9[��ट ���	�5�<�a)����I��X�¶�zb�����?�!�KM߼hd-u�����yd}�~;�?�'��(#:w�kE�e�&h��VE�8/��{��+/�GIo4x��^����)N���=���C�d������s�'�zQ�N��nx���?��?�|M`�1o�W�2�\�cm<��6:�+�� �O�/�:��������6Id'��XZ�PT��oB�9S�z����������x�W��4�@���i��AfVV��l)���$�� |���?���⧀��C���~����Mzk���ud|ߌ�X���4j����+��ٞa�x�g���<#���[^�Vk�{��p�_��H\�c�ɮ���7�6��B��dZv�����y#���j��WR��plc�z���jW��l<m���R���t���>�iZc!>ᇾk�?f����ŕ�eǎ��C�k$�LU��e����Oƺ��#9c*�ʕ���O�GᏃ��S@��_���\�is*ݕ�?�1��kO�D0�WWX��b@�H�($@��=FGǯ��u������\�>�چ���"N���Rn���>�zҥ7�9�f_�������B�R����ܠ��G��a�{�?��H�_��s^uO��<T��2P��c���q��!��y�=G<`�t��4;d��"�FG�z~-��jR��K#�`�����V�?�|��uћL�������Wn��g֮Hʶ7�������R���o�??�%$c:��� ���^� Z���E_�.���0� �R��^� Z����'� r��-QT{AMju5�}+�?�Ry�OZ����y��.��|��e�G�omf2~��Î|�i˲81�S�RZ]J|�6�o���}�nb�^Z��>�?P�7���^���1#��[�����=�[��RY{z}kЯ<;co��#�S��rqԞ��.�a�a�օn^K�M&�����|_�Nx�>�>��G�O=�$��r��|��mf��ҁ?v�^��g��J�9�n�����^��H���d��\�.�����qU*t1MR��[���b�����f�H��(��qޢ�s�q�Ƭ*��� k��[�&���<g�6>�W"�!���D��?�3W�J��� �eቯ�NՂMy/�=İ$�;�{�qӏj��w���2:TW�l��.��B��cQ�J�cG���8Nǹ~�:���ږ��Kv�k#<IC�v��9���A�7�x�-v��au3*Gd����9#���t�
�%^|1�� �--#�y"��Y'�#��^�}�O�H����	�0���1IМ�dw�MUJTq�WB��{�}�O��s��0G��U:^�TlX?��y���?�'�`���C/��U�Ы6kݴ� �B�Q_'M��T �qs'$��<t�b���v���^	�}�S��1;Z�6	R5)�3��f���]
�FxU��
�$��C�0� ^��S�VZoĻmFs�{i"��#,.q��}1'�Y)��G��������7�gP"��/����38;
�k�Th�7&����a��������f-���V�J�N����;��ߵ���G�_J�J�#���Hbv�e gһ��������=p��H�Ip9©>���~��G�σ<7�#ȑ�2}2��.ˣS�.g�ϼ�}Z�d�G�C	��K���?�+�A�z�Z���z�@r�潛�_�G�<s�Ia`�^��������p�pF8l��ڼq#M�C�w���cUUK��~s�b�^p��K���H�o���jp��'�m�D���.}<��V'�k!���d_$�������s����p|���>*c���F�vҩ7�N�*��N�f�U�o�1����}�S��fp��� �����:φ��WP�� �K4M��[�gYq��S�θ�xU�.�-�3[���jIs)��
 '<�O.��X����'S߹e�u���7�� *��N�NۜQ���u�����|C�������j-z&�۶0�m��/�K�{��&����.�<|�V����\��4P�-��|T���vφ,%p@��>�ӭ���e=���؅� �5"I�H���K�FI��5�T\�cӍ�Яy� ����:m�Ԯb�S��@ϵ=/a��WC-���Y6��I���$��[��ǧ(���H3$��{����hT�1�[�-]*���1��ǐ��5���ܿ����}����%V�[���$5f{G�W;��C7(b���nQ�H'��ɍh@V?�o�A�6�G{~��(��m�aai6V���(θz��;����� 
�<�����s�nz&��e��hv|�S��خ���.�����	Oe������1���}3˳�}`}|���s�	�s�p��56�� �F&B�♩M����W�YY�}S_W,����vDʾ�~r�J*�A���G6�~CwR_~�i1�p�a�#�_*�����x�;��P,"�s�E�����i��	^��n�0�x7W"Oe�#�wr0��V
�Qb[�ãk���;)3��?��w;7mJ޾�}���6��jс�u�emwK���w�qԔ;F��oT_��K�h%=�oL4V짹T)w^G��§�B���[_��{��ǡ��p�W��r0\���u�O!��e�'�Ո������ R���������{}-5�>���Z*�z[5ے�א̺?bq[Jq�A�?������O�Ѩ����b��m�"�_[��T>�c(#��b�BMƼ_�w��͌`�5��˯�tر���$�D~�L*�߻��h�M;�s��u�=��YLX����/�FzÜXs�u@U)j;�5��#`
ҏ�a8�w�!�i�$���Ǭ��uolrߵ{��@8��*���c�Yh��[�ZH�&B��y���a���,���3��
��NQդu���pf���}��M��}��J=d��6���[q!K���g�l�� ���<�gX�k�sZ+��p�l�Ȓ��
W%�^�t���"D7�,K+���ƪ�F6r��BS���j载��}�f�B�t'f|i�A�sƥxɳ�d�4;wȠE\M��ms*5]��xcP�Li�~�#��<ڔ!D��� `��6T�;�d��	���BV��u�	�}R,�9����)6�w����JL9tx^��P2!�]�5�a�`}�����Rl�%��3�/���<�2ܨZ7|\��Ɖ�����T�{(U,
='O���0Ɩ�^���L+K����A��4u&�����8��v��L��Q/xn�^��y��۾�]�3?̱��"��KO���R���!{�s\U���H)T]�}��8��������b�E��K'��:r��U��B�)���t2W"[���©9�-Z����D�9VlW�7��~���&���B�q�T����\�mw)6��4��,>�_�1�/�5sA�-���k��}o-�Hv��9q:a��Zm��x�/5	��yv�k�nT.a��oȏ�f����|��b[$ɯ�
'K�(|`m4�JrTMY��	Ee��4��-0�ɔ�8�#�
���\ϩ��}3���S�	�k����4����w�,��>�)��1�q{���4�[��O̸�W}����z{R��n��^�P����KIp����_�.��2c�A�Z���l��������`V���+/�����p�Q��՞���D�����-S��uW�`�?^��� <df�?��ƫq���ZN��ڕgR{�=����L;��ζ��wZCG�ؗSV�����P{f1k�U�T�R|y{�rHK��1��Z�З�(ig%��&�;�=��v$Cm�_����/>O:h-��A�r��m���C'�)dg~ܤ�����S���I�������HCBnz��\�?���W�E�
��=�^�nhc`7�k�K��Udb����z������e:V0SVZi�&�de���h��R����ޱ0N�/"8Θ@��Q��x8)��X�[����%��2b����e�`Kv�@�Φ)^w~7�C������"F�Q��� 5!���9�nW�˓YL���w,��4*�k2Ẃ��n�ĕ��j�9��ֽ��J��c�~�N`�M��=��5Q񃵩��\a�fu�ȝ�jY��A�"��G/�{}DD�V�!Y���K�h������12,���ڻ���	N}����%�A/��u|\�����
�n$�L5È���Ϣ�4a7���p�j�w������}rz(�}���pM8
�̒(1!���?�ss �K�!ohq�^�J��>��͎��F�֝���cQt�N?W5V�/�����A�^��� b�/k��̧4H ���v>�F ���ݮ��F�+�p�>�Q�����˜|΀ُ�
�4%�,�%��M�Fd_�8EKCڟF؈��>�(�������?Mv��R��|;�����L����@`��M��i�x�Ce-�N��p��^a̞��8.Ϻ�[�.}{h�P����@`j�0o �ĮNtV�z�Q���o�L�M9/�e����;ӇL������E��G����G�p˃i �%VW:�5'�\t%$>]$3)��9�H]kAK�n��צ��ۻ�jB��ߎ�����=9▄��y����tƒM�B��#[X�v���R߸�Yr�t�����ze�n� OV��}�:�*K�~nw�*M���}����0J���c�x�\<H��9I;�=6׮b�/�"Z}�����T!�N!s5Q�ӊ�Z�j7@���S�,�d�Gge#6C&��J�*1bc�#���ܲa��n���١�/o���<�M��X����]�g�%��7���<�&\��v50;�o?<�>�?Xm��g6�>o{�'Պ�.#Z� �1����/��Na%��L�\�^�bz�"d��O����~@(��L6�:i�4���(��fr�d{����ow.���80�A��M1�Ŗۏ�w�'�u��7#ǯ��M������M��t+� ��hd������OD�k�S�3��E�]�-5i�:[�B��.���ߤ%�%�F��"0Qw��(�.(�E�W,�������44�[�Oq� �� �Lqd}B�BQ��͇�Ͱѯ����T
��d�'�k���A��ћ,�g|�Op+_=\*�{4�+|ո(��&�UA<	"�������О>t )�;K��7V�����$�]u���C#��q�����'z��g��[M���I�$_����G(3~ �����e��*��S���]y�����3�~-��	�3��,\\)Gƒ�'��'4�⟰X��ک��1%m�76xE�~x}gJ��Q��hr��~�	�;~N�
N�����x6|r~l��ӣC�(�rW�9� iI��x��,I���o�x��L�Y}��M(æ�� 1���~��1�9S:�P�|�W|3��bZ�0$D�H4,_8�)l�6j�F9�ٳ���ߧC�!V����� :Ro���FKN,�{�G��3����B�S��d[�]���=,�6;�|�tw�N!h�)km��3O2 ���h��Uo�}�ϗWe�\'��6�V��(Zr��4.K�c ���b�J��-��aǁF�������[�=�ɳi�����9j%����N��H��ڴ�����T�!{{�q��h�[�����cɶ<����OִC7��{�C܂T���5�3�eڀ���� �V ��˯�(��YD�?1V��	�߶�УN1�{]������������Gg@��y�'A��X�h��b���T������D|ݢ�5�s9�Ho�k�����lڃ
r�&� T`~�+��M�v:��L#������q=������.zX��������,������}���|��M��[S����8Z�a,��y�]�-RG�^����υ�[�]8A���݌=k�J������B��&X��Hr���2-�����Ǐ<\^�5�&�i���H���W�'�LM	�K�����ѱ��Iu�2uK���`�^��N�[X�Pz�z�
B۸�vt����n��eB��s�^6p��t,kL[���N�.�)��~�.�	��;�N��M o���)x�� T=�W�.�}�n�;������2�U^0�2��c�B~�s��i��#j'�KNhi,ͭm���mLmH~����e 3
�����a�@D3-Z6y6t���y$���?��5��hH �W���{�@6���@�s��eܫj�O���@'D�^�W:	�V��j8����A ���L��_�zڙ5%��'|��2G�t9{cӶ��cU��/�45����%� �Vp�>��_ؗ�z8z�Jծ����>(�3`������Ut��U�ef���-�O
>���Hh�.��s���*nE�0V%ۯ)�6y��z��
�x��vk�0��X��1֙b`�hZ4�ܕ#+���{ �N���[�N��!�V	��c+��x���}�h�a}�^8O������9*S䔌��_�(Z���|�ŧ�G��j)�t������>�f:K�#F��6M����JVP_qw`w��9�z��	�0f��<�X���o���D�S6�,�B���2���o*����
rJ���Kg�wН�c���ˌ컾��~,Z4=��Ȕ��))������*������7���k,���d{h���otz�åJV�m��T�t�Q�e�j�g�pd�|O�}���^��F��dϯ��I��ʛ=G`��Ys�ɚ���k���(Y�V�G��@�A��Eƶ��v�M�_rd6�������;=E�D��1����A.�&R�l1Y{�M��.p�{&���*�T�(�!��+���%��0���Mk����?�Ltv��h�l�_:�o�(�N��X;�#��-@�ٸ� �P��iD"��qhdKf���]���ؗw������
�>�si��(Y�
G����g��o�P�%z�De����Ty�̗�e�2���;݋j?��E�0�CG��ul�}�|�vRNi���D��YnZ	����.Y��3��7��#9(su�I����Bm�ET:�c���J%6f���z�"�TF��*���~���N�IÃ2�F7�L�P:��돜�.��-@hU�s5�d��fR��LRsrh���U�e�<z5����c����z�@.Y�k<�!�>K��X����Y~�p����:���8r(����)3%����0;�5��¢c��e�"���b���"��Ϸ]�N��k���h���Ɣ��1߉t*��I�SoG��!�{N�ؽ��]#�޹�����n�NFY��I��!�S7W?������f�ѣ���>-�mQ1\l������IwX�G����ґHw�^���#�B��o�k�fX-�y�M��U�$^r}��.�KkF�v��>q��x��74���!֣�}���Ѓ�/�o3qW�E��Oa��e�7"%[_j��2�aŻ�e����ܺa�z����	9uuUʕ����]y���u���)����l�tsZ�c���NXL��۟��/�Pj��~�n���Fub�o4y�3�U��/�79�
�ݒ�bB������ p�6�08�����z~�*Pu;{�q���o)L��Iu�N����ʹ;VZ�W
K�1]�Iϑ������?�>��:M���8|���tc�+��Wc�6�Tg�.��n䲵���4N��?�N_\���S���� `�?��F!?w�t�E@�d!P@�V���(V�FaZFfS����{rL�?�
���'#`�sm#�Z�h�J=O�u�|��ƞ��O���r�N��n�W{�fZ����c��<���߉gC"��#B�� ���s>5�x�$�jQ�?�h�I�]f[������H�&���z��͋&� �	��at2�I�K�itk��P�֐�T���&c�s�d���?)�a������iݴ8���*�-Q_?+��Ȍ�4#!�+2��MψC�g�X�F����&Y�涴9��j���5k���z��֪hٚ��Ŷ`V�0)�ؾ_�����4���2I�Z���OC�������kl��J���L�n1��5�n�H,ޝ�~R�F���(��(5Uɻʕ���jx�Yq�����	�=��"�B�r����sw㬘���o�Qi��$��̊B�{k��ZTʗՊ�����C�� ��+���
�v���tŧN�ȣW6�.�"��n�|�A���!{z�|ERo	� ����_�e�*"G�>4�}��!��"�}����9tb�zn(O꒻T ��>Y ��q-� �
`ɼ���jRzE3�i�Y�gJ�K���}��.G��׍�Nݵ�n;lZ��w�Ҟ0K�oU��@�< Y����1�a��~�?2@1~�qú����C�������ӢJ�E��ޫt����samP��"{���8�b�YC��t\'�k>�ǵ)��Š�. ^��5��ҟ�����׽?��L;��������$���{�c.��m���jr�9�r��zÒ
lm�R�Ųb�RwRp~E���rNm��+��/�t�����7�B��+z����a-��k�&L�s^�z����o�&0�A(Z�����٭Rx�c�B���t�D�VЍ�9������T�!�߶�&�� �JQr��Ѥ��W���_f8��v�d����cj7��T���<��ta�[H��ܣ�C�6���E��K�s�Q�'e�>JX9�e7]��<R!w�b.�Q�~l�.�����g@��;Vhlt�>�n ���_$m�^s֐��dzfԅ����K�=MHO�fo���j��iv"�Vm`?��ݦ�GWk���B[�P��~_�l7C@1���T\�?�cjT��>�r��4?�P�^��T���M;t1\�R��+x��)Q,�G�J^����fq����Y3��H�d`�4�E[V2%�Q"C����U���M��\�ד����sZ>�!�H݄�����;�o,ݹK��YK���b��i&�5���w_s�c�t��;���J�rvƽ�V-�w�u�f���|��x:ϢFB�L�Kҵy4�F��v�iA���L�fu�Xɲ7�_oﳢ��gIѴ���,��dr�ߪ����H2oJ��S�Xt-`�:�Zmtb�;mݡd��B)��I�$���׬P��|�����%۸(�p	]h�j_��I��7g!:ߏ~Кy��R<,�$�
��bH�~�n�]\*/W��D�﯅�i�Z���_�d[Unyʓ^�ج�,t��)��605;��3���U�u�$�h��?�a&�|H*��]���x�l�׺X�"�p��P<ʍ�����T�S�]A���(�g���,�!3�mx�p7x�- +���x��m��U5w�*M �_��'��!�������������x�ԉ!��֭%�@���*��j���T��V[��.S�~�LT���e+9B'��9�A��T�x�q��۽~��V����~��߆Z�I4�	�)��t�����ޥ��b�4g9�j2�ÍvS�^�{<t&@�l��k��x��~�����7^��U'y�l��Zz��E�r���nUM�?��=#�`�:�����Y�V���������PB�`Þz�$�{ �X�8�S����= ��j�Pg��WmB�g��}b�s;y̒�A�~��`{ݵ���:��|�dk�"��.|����L����1��7vNѵ���0����]��!\З��;��1V���e_2�p������1�A�4��q����l�g�쏸�Z�!C��V�Aq������Z���W(��>��	�bnΈ��̫�	�m��9�↨���oŕt?��n{��׮1(�#� �qB	�py.���#���ǧ+A�����;QˇcQ7�e���Z��d����d�
�R���t�TdlP�%<=��Jw���r����L�?��ʅ�ֺ�C:_��ު=�@"dl�қ���}��KtLڽ[vU�S��a�d�r U}����������Rw�����CD�/��C�a3���=�)��{F�)8���`�������*�}e6��fQ�RN󌐾���e�4ݹ�Z�R����z�����T}2�նFl��剴����_�$�#�^4q� }n2I�|Vޮ#^6���$�%r$�De��MM����h%�B�a�����ϥ��'�f[v��V�!#&2X��[|��W`�o�ԖbS�}�O!�[ ,�o���RtWu���~�!wYp���̱V��l�<kR�3sa���NE;�)y�RC?X���_qj"5v���z��\0GFj��޾��@�IPH:R��ުHb��k���ث`���`%ʀ�¯
7+�rb� PZ�QV��yԿ�TLM
���O@��t��Vա�bM���e'*���
�̧��z�5��n�H��ꕑC�fV�,�����U�X�cs��ݖ�hy��6c�V�'���{Z5��Oi���Mm݀
�������fۭ���`B،��G�E��̄p��Me���d�<��lO�+�T5#q
�0y�W�c^�\ϵ�{�є�I.T?$��?g����3����r=f���X�2a�~y#�6*�0_�1c2 ����#l�s�Ѫ�c�k�H�/���g�ܘ+㯮�����T�E�#���!�;CԘ���)�:0�Ny�7C0����ƅN�͑��D�앛y�+e�3M�팇����ͬ�
$;5���,�vg�+"��fS��c�?��4╥#����B�?ǿ���8}��1��?Oe�9u/��6����(mg̀��ߘ��	w�.P����e�,Y�-�*��7���MW��[�_c��)�k��m���C�𧢮+�rT�5��8���Ӷ���cɥ,l)jtr1(46����w�U�
 ��Ѳ�"�=΍��%_ �<�����/�X��,�鿘�>u���n�k�%|ez��\ �Q�1�<�o `=����:o�f��J��BN,9?d/�|�{V�`#��2�\Mv�iݴ�j��i츜��Ʋ�Äx�w�v�:�ն��xztd��:<�K7+R�L)�@~+�7d>���[%y��=�ϲ�j+Nl��᩟�!���aW��x���(��J�q�ܥ��]�����{�'�P������Y?�jh��\�OMJ�i�cHK1�w2O��֛���<�(�u
���"���L�g�@�$�$��Dɪ�d1�q/���������$N�m�.Sq&�VtZ�r����C���5�u�&����9�2}�wd�3RN��zk���sT�i�����}��͑W�(���OT�����z����ް�Z$-�gQ#��R�H{�s�Z��I/�W��~r�������I$.xX��v�l�o�U$NH����}�2�Q�T��+b��*j\�ħ��j�?��b�+�Z ��5�yy���E	E��=�5�ƣ@hX␣��SRЎ̗v�ax$���Σr�,��o� ��f��¨�6�S�J�B�б!� �ҢkMJWt
������ _���֚���]ݵ�d����#8r衼��?pg�k'>�b�\@E���&��UH	�����}��dH_�-NZ�ٝ�;ծ�\L���B��q�b���)-�\:��y=�7�7)��p���!�U���F��&��Uk\j�2b9l���Brem��\@@1�}/0��~�}������@T��_ZS=~�bs{���-B�
87���9َ��3E%�W�Fz-u[7@���=��ޯ��ԧ4��h�D��!�(=s�Ɗ3>���	����pQP,���/�dI����fs�5�����q6����;�g�j0�Wh0rabNg�����O����)=1�B�cV�>(%�&��Wq��%F'+�ckV7N�����^��7�n=4�0KHҁg���ʅg����7<^�]w�52 K��C�"w� �呂������6@��;���T�VKY�)�gp�����s�	��4�h����=�6��u�6q|vX�8���f-�k���з�Z�EGCK�vt9�����dAX��3�W�I�>u�UF��w9@�kΪ��7SE&,�jO�[��f�K�Mأ4�{��ﳜ�0\�W�do���|�I;�=wi��
��c�y�;S����]`N�4Q�hy��$L�6�ae���;M��Df;�\�s�-���c6آ�ӓRc1Tk�N�����!v}���tv�B�R/��'c�w����	x��
���%�w
�2�K�)�ddo���Y�!7���ֽ�3���zY�j��Qeԧ��"�	�)"���`w�mXv@�A�(�ր7u����"7�W�����?�=[A�9��8��E<���Ψ�%ҹ�ҫ�Ɩ�'}����>d�2�ΟhnJ�����)�[혞X�=�3u�����7/u��BeA!-�
wI|�/���?���aoj. �ze�MNV�����aE�������:�B1?�WЀK��P��ʨ2G�Q�PYP�[����/�%�8��C0p�r3P)�;I�WTJ4��e�8$��Q_�P�&���!� X�ĶY�;����#ς�F�S�6�ߪ}��1X}b�8/Z�~+��K ����
�@	\k��t�A��ܚ�^�|�/s��1�yQ�q�ܷE�9[U���^�K0����]�1>���j(�8�3M�ӷ&P�R��1&�f���B�v���`��x��jw��o��)
�|i��-`z�Z����|<-�9��h�'����E��1]1��1����&���<IJt9�2��-s5$T�G����<�vw��]�i"F�0��V�p�'��:6�{�]�!���>� �k��/��J�K�~�"3���H��u��&�{��`��u��d�~�RV��o�|��sjk��W�¥���2�$i�C�X��ܿv�J_��	ք��#ͱ`ӊ�6���:j��(cH��r^f�1N7%v��$S(����#��O���L��m�m�]0���KjC���C��6]E������e�b.q�F�\�5�.��`���N!�h2ճ����d'�1�'�^k������~P�H&!7��b���TV˸�����Z��Z��������Fv���ҝ��3(����2ˁq�b�[Y��Ȑ�3��B�ҕKBA��M.#��J�1y�9�,�6�_���醝��O�s0�䔕r��4��W�'u@8e���8r��<�^�I2
��(��h�J�}��R}���t]<�Lz�<W�J�^*3C�>�*㻞(�2#����E��)��ڟ?g����`>�lL�A���̀�TU��12s�OS#�Lg����G�m��&��-��o�MpWyiH���$q �-�N�Х��x��/��o��ʳ�SV^�3�s����|�n���}%y٣z���g�~y�G�S�{����e���XV�_���H�/<0��*�64���R���������\ A9��sS=Cej��2q��g����|�����_�=��'_�c�X%��*/��w��Ƃ��l�t��/
�sz�;��b%ipnM��9��z0:ݺ��¹���D��L������J�DyUCݕ�h��i
:�'T�]7�O�����Ō��L�(V��n�]6��FP,1&�?ϑc"5�qT��v]:SVҿ����1��&4k����{@�*?Ԗ`��,h���G�i�i������E�dn]�Lݯ����	�&�����/"�V��Ca���/�w��i-��r�z!��ˍk)Q����<��f������5˿��2���Pnl�:���@?d0�q�VUګں�:-�G��OI,-o���as6���$�O���x�mKT��p�诫�g���o�w�����Cj1T�k(�Ln��V��Ӫ6�{�QF��̖�{P�ϳ�� k���D:��p���GH��Dh-=�%��5jڳm�#����c~���'����v�c�ơ=������?#YǷ���?6~Q�yQU�~�Vʵ��R�|���64hI�w��[	��[��J�A��V��>���ZË����0]�Hb����>I��{ ��	M�܍GKҞa��G���:�]�i6�>����*~&�XS�P������·��x G�=)L�hKn&�[Sk�Xt�l�Q�%�3�� �y�(!CL�5^j���?�����=U�~�!_�d9i��0vL]DPa"����R`+٧����B̢|`�4�q���E�j-0��Z&��a��Z'����3�$�!�j��m�*��b�ds55����j���xED�|t������_?�r�[�!����d1�E��XxXa�}Yl���4�&C�cRN$���o�g���]PCW�b�����vG�bx3�D��+������X�������[��}Mُof}Y�7e��
3-�ț�S��ZYѷ�!�D,ŴCc|�h��/N�R�-�i��R�ӛsEͧm�#���?�8��v�jAx�d↷X#���{��钵w~h��s��kXU�ޒf�yX���2c}N!7���&ׁ+�IU��hv�t��iB뉬$�*_z.���L�F�Yw �MQ�BL��}o�M0�3�&�wB�)�W��|�Q�.}L����ǇHvY�HX��ѧǏ:hn��?�^�zf�)�g�uC�eZ�:뻟��
N��Ⓔ{ "Lq�]��
+���p7�J��[%ӳ�_�-��9�O�e��Z�86��s22�T,�ɋ�m�4%��i��?a���Կ=�X+���� z�8�8������:*��zV�pua��Gh�Ҕ��t�J��Av��N;d�B8~���\�$��u�����f������1�uy�ϊV9��}�U�ȟ���(Y�1Ձ�ӳJ�c�l��%����7���(�8�1�ao��XR�/z�p�G������\���,\�^�d�.����,��|�`�����-gk����k���U��[��'Z�ѡ.�m��S�]���؝�5�����󫬭�E��^���J�2è:�=wA%,���q���bc�����aA�zo ��8Pk�%x+�(��F*��ԟx.��(�ҕ��Tc���E��[/�2���9��\��v8x׬�62D�ਟ���M>������F$��A0>G����!T[	�ؼ���>̌Q�Rl���f��k������pݓ�����/O���pG�[�e� cy��l�%��+���g䀘hĞ�ǥl�ȅl3ܐ�An ��Bv��z�湑ȧ��A>�V_����)m<�i����˦�L��JɝPw<�ե�y��}�Ԣ�#��'5���6��⍍*�\��(%�������X7]�XU�c��1\n��HM�DൟT8,�Xw'."��<#\?G/ΩTc �1!R��~��R���Q	NmB���)\L�Q�Pw@��V&z�N���;��Z�� .���8�'I
ͽe��
�`��8�����tN6Z�/�W��ı>�D�Y�3���^�-�O6C�ti�W����ݓ���Ի"U����	|972�;Ր1@�%Ϩ/�YZR�l���8�����?bT�}w�~t���ˆ|uiAo"��r���缾U.}z�g��ؕpx��L�y �چ2�F�.�f�p�W��q�������9D��y�ӋZ�,�5m��P�1�j�������+�2y��b����,N�����2�;�,vZ�~Vрcp?}2UK5��Qy�`|��M!��8��p�q��� �fج����"�&b������0ǋ.*��P����+�iM��Ĥݯ�����
Z?{�f}4S"�A�@�����2�Ѻ}S�a3�5�ԓ)�S}�Ii�K��4��Lt��1��7����C������Ϗ6j������Uwî��Y�n}0yk�@����A=��_�X��~�Ꙡ��sc,��^���ņb�.��E��违q�Y�?�#)�,�����%vY)���~���}+��{����%k+��\�G����uR���jnh���h�#�����/���%f>��(Xl���aFT���*W8L�= *��� ��"�N��*����\V��&��P\�C3�}*@��Q���Gvy�82l�˳��D��~�	�?f�H�;��i�qi��=��By$ �*Hl)4�0�E���R���'�,�/�1�^�r�*��Ђ�}�~�,4����|���-�-���w۟ܪ��~�K=�`�
녖4�{���.��ݒ��>�b����č�(�@���X��R�t�(��/=�2���^�}�4LH؇��͸�{B�T$�.�))��ze(0{RL�y��z\>Zf��i�/�s��L?��c+1��ް�"s>_�߃��ʾOI�_@6ɞ���ʝq&��9T=���L2���2�%2��G�_Nc����l��W��ۑ�Q�=�;��%�hƥ.$nq��a���O�HF���9:;I`��IQ�f$'�t�ґ�me^/�lJly������ƗT;���Vu7� #��F0��=wl���jQ��!t#�o�Hl�1���_vg�]@-�m	J������k����֨���^��J̈́�B�sfZ��IG����O����;�ʼ�xvJ=��Ύ�Ceظ"�v� $-:?=??�3�:Ւ>��j��-- E�o�:�QN��v���Zkmw1*/�GkW��Avs���!�Ō�2k��˭ְ�� -��|�>���H1�T��ƺ�����x�c�6޴�>Ӛ��5x���-���b�k2bE�wJ��csen
�F��	N��j%��T`�cz_ile�]g��4�zUmd�[7A3��1F�#l��kK�i(�����t.���Y�<�D��3$.�����_$�qF���$�8�]����uE���_�
��P�.����H��H���y��b���S��?�z�ڢ��7�y��u������ա����d,��j�/�����Y�r���~�C̶4� �*k�Z�1�؄7�f�� "3�rd�	G�9�P�,��V�f�1�cpQ3mMä�fl�8����&�d
w1	Ϟe��\�Q�*�9R���`���v0"���nJ��[J2�~m�
{�_�C�Ug�Y����(���`�=6���h^Q2�Zջt���'q��U-C��k�@�`�\�R���9ya�x�~h�w��k��o{�����z��
�j�lL�:�!A	W�~��шW�#ل,^�ݗmU���:[R�~헵�@.�����i�G��y���� ˪	�e���OU��D��I0��mR��6���5
��>�ze~q�pǇ1+�^�?���@��;��9�f+���G�Gq27k!]k���тK�By��E�
��?Z��/
z4�x���� ��I�L\�|gb�����IQqIo\�^��ɠ����>�)�i��M���G"���hO��y[4��j��O���G�3M����M~�!uk+"��z���h��xO}��mIss޹N����K��R�y�6�yg��'}ʟM|1�E���ᒹ�:�h�����{������Ŕ�ꪰf��ԃ�Qi}3u,4n��%(��O @k������;+l��)}�I�[���Pk��JJ2�M{�w��w�� i�
��7�5e���am���$�I��Lq���_E�I)
M�oGUO��ٜ"N�ąl�/���{���ؘ���e�r���6�7�rci�s�hyZ�w��|:�9�o�4�X��m������ 	N����^���ӿ�ZW��au
�'�Q���o<�������l�n,�擧Ҫ�H�Gǔ��ݢ���^
5r(��,�t�⻶��H�����[���*�P��������O�`,��9lC�n���qF��kNʤV�!,�m�r�D#S���yc;�a�ft*'Mz�ˁ/�GQ�sq�[��̶,�V�bȵ ���]��ʆ:��*d\2<n�<�����t"+�������n��Q�
����%���������۸/��89���ߝ�������GY)�i�"�'�Y�?j���k��MF���.�YW 	�~ן�}B���7(���G�Q�XEhy�)�
_]Whŭ�eU�ʯoM��릏��ƺwr[���0e>�Pd���|��v6#���I	�c7]Y�,>���I��ڶ��i�`�g7�� (��>�E�ȵ{���́�R�b�̺�dt����Ժ����83r�9"`ZLÆ|д;X�g����9�>���r��-���6��8a�͡�{�s�GI=�G-r�Y�:������r̿�p��W5�.����W�C¿$�NZ��(Q� :,?8"�/�F����L�:���2�$�򐁼YR���t�=����\F�@�=89:Q#ܠ@P�Wv�BoN����`�6B�8D���x�A�j��U�]����W�t����Y��G������
mW�'jiEZZ�U�����\@���!��J�"���_��~d��c�ƫ?�t�֗?�4�|�}�����$e!X�kv,{W�|��&��~+k�����.� ��'	o�ğo�ϕ|B��7��M5i�-?J�>f���v�� ���߲�i^$�g��jZ�vj��e�dT�"��1��*�u#*�(��p��U���fd�w����� �g�d�Ǔ[�%��|<��#�0Ijۛ�p>n�s���hi��'w�|O�K���	ޯh��m��6c����EP� ��߇㴒���g��K�0A� 4ps�9����C�([x|W�?x�[{f�\����؜���`O�@l�l��s�c��Nɭ=Q�׆�9A�/�F�W�v��hw�s�q�͂�9���XI��I�6
�~|l�4� x~mj��/{���tY�2�)?9R˗=�OL��_�|<�kk���0[F�\i���g�O˸�;F1��޽�����>MSG����7!�G.��2DC���|�y�EDq%.^P�kz����:�������:G�I��h���Q�V�!�d�`s���צ|7���(%�Zu�7��Ix�wIH$c'֭��wG��݆�� !���ؖv1B���.������+���&�[�O���V~=]U��Ks�R��1�Cv��ڶ圚m�q5qJKC���	U�?�Fp�5�����Y� 5�/K�ծ�t-ᾈG�2��9��3^��s����{ƞ!��5�d��ɂ�%*N_����ן��çƚ|:���[ߟ�E<�;.x݌`��\�$��h~s���.r$���9^�[�u)}�$���E;��89�|9�,�,����ڼ����s67M�1g?'��ɯ�?��x<?�3�+���$al�A��sֳ�,h��U���f>�s39f����2��x�k����NX�� kY�A�Eb��؃�?���"��9�b��ú]��|���ݹ,G�*�.��ץ`�����+�Fz�[<>1�� ��$��J���Z���^��������6��(�c��g�d�'�&u� v:�5k�?�g���q���M� �G_F/J���?y�ܩ�EU��S{ө��0��� �ƾ(����ȴ=� ��� �޾�n�ھ)��2�,�c��� �$�\F���Y� ���G����r
/�֌o!�rv�3�ڴ�G�t�;{
�ۺ_�_;]4~gR-h�� ���
as�Ӝ���f3ژ�l�:д��Úc��+�u���H�� �>�� ��8�����sҥ�۹5�j� �=��nG��5$���Wn�;���z�U��e�\���ZBaֵ�au���<��[#vPv�J��� �Kl>#n6���A�Ȯ?�B��5ӒH���U���{�W���5�a�x[�?P����`��kN'��\��>�+ʫ����[���C�3A,��(�eS���?=F��s��.������^��m6�C���S��w�1���·�v�q�}�#娓�=�X�O��D���}8�(f�H�nV{���3���g���֝��ZO�'�4��.�Y�����u�:��rMj����A�e8�Z����;�_6���_ſ�V���Q���1xWf�|�}��������`�g��>i><�:�Y��W�����7ď4j^����TZ`��'��~�et����/q9�|� �Z����x(�j�z�@��+���18
�~��~�����wM�K�3��'x.�q���؎v؂}��~-x=T���lPHŷ8V�K�G����Ǝ� g��{ �$��0${�y�����L�}�3������/�s<���تp�7�ϙw<?�����L�^�2�a���K�$q�~�$��I�p�.��u�֬���il�T�rE�!C�}p{O�U�)���ה�~U�IF>�Pٟ��R��Q+Ǳ�xWŚo��K�V�lS:Z�.F�c4���|Y}��ٕl� fѠb@� �`�3��	-�bn���x7�����>�SӵD�����R����_A(*��sħ^�=펆?�z��5ɣ����_mm�h呎21�y�O�oP𔩭x�xn��L6�ynd�y�G<W-�?\��Z��+X죄y6q�I
�@�%�I���=>��ޛ�a/|]t���,],��	�~��y���o���j����ռY�.-��%��j(�}"��&��c��V�������7�>+���/�K�i�����}'A��Cƞ2v���c%��;����^�z}+K>(���[��59�mc�^\�� ��v���Nֺ:�)Ar˩�ͤ�k���d��܀�N1��U�����1�u�G��=g�� ����f���j�d�!+	U��~��� 	��ٙ�5��p՟򫊩mPrB:)\�GՌaW���Gr5�Ƙ4�c���}� �ޓ��\�~:�m��/�����~�ԉ㿆�d/�|�vWY�?�W,��rA�:������ ½�w)1k��\}k�m�WR�'����]����3��^��� ���q�2G�� �<�]d����l��C�]��iu��h�2N��Fq�û S����iB�S����_;Y,_�!`~ѭ\�;I�S
:~?Z}����!��ĥI�bkS�Ď�s�OLs\��.o�-$�H/����;�#��䚟K�����9U��x���k}p0<�g'������;9)ݵ!��~�����~)(����6��p�z���� Zluo��?^z�\��N[H�vm��q��7a�&�Z����.��� �� ��������]kE�#�����L�դ-��'��H�>�&��x���>����Վ&�7r$?�d���� �M���ھգ@8S�1�Oޖ�K�?:�t�[b��&����q��X�E��û7Z��Ij�����y�#L��rs��\�%�a oj�1��L�XѼ_�	.�������`�[=���2T:�~\�'��O�q��q��:}J��~����r[k��м;o2�L���Cg����\�W7��̑]�}��C2j f#îz#vǦt^&��-�HV�Qu�R�6��Z�E� �я���.3�N+�m>�P���h�/e��myI꓌f4be�#�O�e'����:߂���Oy�u�.��^9g�g����V��;��� P� ���V�}���V[�� ����TH{ ʏ�j�KV��i�N���kkj�g��6�Č8�\��{�]t��BDK���g|���It�{��<�*ꥈ�5dwQ�18x�q�����?���:��6�^�ӵ��j�RKq��Z��T�ц��k/�ƫ?�k�x�X�&�</���!�K�1*�S�@G��5�ֶ�F���5ԯ�⑼����b�c*��dy�5�2���i�֤�xt�VXm�sl8W�pA?Z�R�f�G�<}i�\�sԾ~ך� �/K��"��F���ʀ|��*U �WI�oۛ[���g�]�q��x�e���IJG^�iܸ�A9��٧�k�7ŏ�� �z�����Ind���
�S����R��#�[��MQwg���x��
8iJ�V���r|���JsI3�>1x����ǔ�30CGh$��w�#|`�6������~�k���b���\j�ڜgv?�����"��?�-Lq������4���t�%�h���#珍����Ə�:��4T���H����	4ڥ�O$dך�'��w����V�����<�,�P�sۃ�k��b����&�"������� f�/�e��km�d� ��� c[�e�Z5�
f��������W�/��R�����F�_��V��c�m��1,p��c���I� ��J�M�:���Ԓ0��G����31����h��*|/�ثY_��?me�e7�����+i��_��~��S� Z(�Rl���|����� l�w�v�4;M�����K$�9ۼ*�^��|�����������3t���w�nX��&	VӃ���ݟ����RTӵ���88��� ko���W��xr�kh��&�a4�R��5��!���MY�.e��x�$��{���j�\�n{��@nc�X���3�l�c�	�2|լ�C�>5,����k]Y��8��%"Ks��;�NT��j��c�ޞ����ű�i_d�\h��n���(��9e9q�1\\�呥�|#�Ճ-嬖yu��� u<׽:�����j�ڵ�j��}�D������ǆg'Q���� 8�+��%��Z���埆��7{�\]�b@� r÷j�t������N��oI|+6,� ���5��x���K�C<�Kѱ�l�t����H�W#�
��&xw������׳��E�Z_$X�.�����$�!ZC����q\���-+����A��MO�X!x\�����fudp;��s�~ X�ipx[��:��s5�����wH�rF}sYVp��T��W�'��'a��J<ԡ�ٽ\J�NX�7<[�o\����;���E����4�U�m�q �ҳ�H��5�[����hKV3��j��8\�
��<H������H_J��o#-�A�z���<Q��i�f�i��ֳ��Vg����P2q�sֺi�kL��NNSf��<1s��]�֛r�2G>���y��K���=j=[�ͭ��;X�V��_��0_���ވ
p�ָo/�q��pay$힟�H!_/n�o�]I�s�x�S�{�>3��c����f���%�;�}˴�C�>��^�&���kW��sj7V����/!q$��Yp�[� g���e�v���D �`c�o��Ts#/���C�"o	��a�xf��WH%y%����݌���`�>�v�_�� ��?A���V�*4m{�@R��Ps�.pq�A�'>p�!vd'���UI�d2����ߖ�Y�*j�v��C�u�Qꥴ�M��$�!�#m��� N��Il㑞��͓wkuq{�L����ѯ�'��?���#���?0T~|H}mt��7��Q�;tL���s�#t��0<1���:ڝFE�)�Z��-���m�br	9�?RN	��)Q�+GҩF�=�6b,rj}�Z>�ܡ�j�����8�	9ʜ�=��U_�r���F���0�8� 9��-������m�?�u{)�o4c��q�����>��izU�jP=�­J�;$H/XH3�v���t1�M���oP�R�W�V�*1��Qvw;��`�U�o�>��|[�W	`����ǯ�v���c��lu56�5ǴY:5���A�W��F}�ޯ�x?E�i�� ��
E4��iVLq�����x�Wj�7�T�އ�|1�S��V��� �>���7E�Οm�K5�l�4*>�j���ÿ�$_kv���k	yv�Ie|ځxd�l��'>�c�c|�W��"|7�ǁ���O�]��|��cv�1ܱ�m
T pO9�:��_��q��6�xR+W���[ym�1�9m�Ǳ�y��{p�j�t���1�O�|)�]B����;�:D�l�z�Z��C;a�.��ז�w�/�4?��ǁ4�d�n��r���r�FP�K��l�rs�I�xk�7��^='��֣���6ҽŮ��¹��`㎻��+O���{ačW_�Z+{����X��KG$���� 8�ڦ�m͙b���"M������� k���\��6:�c�����[I���b�<����~8�+MԬ�"i�����^�ӵY:M�1�������|�9<1�i�ͤ��K����NT�0+�T���>>�T^�L��o�Ss�s�ۏ³ɢ�ٽ��c½�h��T�sT�m�QKg	*xn���^w7��U��H�����P��9@�\�zW58��9���aUZ��W��v:<Z����m6^�o��}rEih��{ϏO��n�d�U�"#�V�W��� �>~«kz�H����sQ7�	� X����$���Q���#=H�'�[	+�un������s��(��(��}5�����J���MS௉t�)o/��QFn�T�.{�'#�޽O�'���|�sV���#���*� �~x
=�'���&$� ��s<#���f��m��Q�|7nluk��������r:��\g�)�
6���aFG7�?��+� �����MQ��ڙ��W��}����.�v��>����h�9���+����G�	$t> ���?�7�q�Q7�_��»���9�=�ѧ��<�@����� -2��~�k��� c_������bd!�$c$� d��u���١T���S�.��G����(Odt;oS��D�	<<�!�X��7,wQ�_�#��������WԷG��3�A�W�/?��y�h�c�hT\FH�#��]8,ʖ6ꔝ�s��2�^Y*���o�� 4c�7��ۓ#��U}w(ܹ�{�I�o�?�RY��5��rs5��K}��I85�{5�������0�'�,���<�}y�\��mj��P��+4�h��C�Ř�l��=?ƾ����{�O�6ۻ����:������p�8��p��\0�*���Nj����5w�D��4�>$���֨|g]�~�G���}sE�q������a|��(��>�'��V[���m&!�d��Y�Q'�4eݷ6�=OJn��ض�uwu���F�d$|�����Ҋq��.cɭ�{���c�Jҵem�� ,[����XPB�f;T �x�j�C�5��ϒ�iRj�p��;3�� �g��o� _�� ���kҾt���� 
d�r��� ���^����G��O��?Ah����
kS� 0�_|�����;�#��i���+����|K�g.߈�G�t���d��#�l�~ v�/Ty�����?(�B�D�����%�C/z�dna6��k��?2�-I�n��OJn����R,��	9\�TR6ن�O=�f<㦐��H�2g�Lm�\��,�32�cT]u�4�p���)�`XpG_�PH�pl��ai�5��{oČI�3�|�� �#_�.��+��aL��?(��?��� ���[c���ƿL|ƛN���>Jq��Ex9Ź��#�N��ȭ2��ʒz����r�3�q�L�h����T�&v�5ޕ�{55c�]�)�$,cǖ�$S'x�$�͒�=;�����AY�F7.�	"�_��4���^�$b��V�� ����QG~qX{
�j�=�s���?���;����� a�v\x�TV���r`s!��q���|�W�:�0�$���0.���z� E���9����	���Z��1�sW��U4�afγ4���.� ǃ�O�}�wb�z%�i��cH�+F(� G�q����Z�qa���^�ݘ�J����s��v-��c��!���rI�:�+���HB�V�s�\� �rz.�[���KAp�E&9u��m����]�+Z�>Q۷p9�x�O�Q4�� w+v?'��|e�	2� h�J����=���$H�� ګ7�^+�|@�� 	v�Pg�&3}�#5�� ��:��`����_����3bo��ߣ<���h�B�H�VF�$�B�A�I�`TP���G�%fX� �� ��J�-I�~
h��^"���h�i�)��y�$��{uv�z���h�>��"wzDͷ{/��O�,P^���?�B�x�\u��������6�ƞ3{ut�m��!�]I�����W�=
%���'��Yc�_>����v
��S��ҹ��SP�����L7j�DV�($��!}�Z�]f��Ex�j1��Ԏ��Z���˛��H���ԇl6���^��I��.���?��Țm�VU�%�t,���Ԟ0�4�v��l,�\ND�t7�����`q�ҷ�;��<������A�\wR@;W�ܒ���j��Z��G�>�|/��7vv���� ��ws�>��}�î��Î2m���Tw7��PB�<|����I$!I���g'��ס��+����ƍ��,	�����B����˃�����9�b�����q��+$��t�W'��̏���k��\ط9� P��;on9��� �Z�r�#�'�J#�_1��{�|������T��[�nY�����[�?�C>��մ-?�n��럯NV��dn@b���¶/�je�O��u ��9��*y\�L�x��^����
xf����dT� ��mW|�3��}}������v�y�\l�<7n�=���9���y������ <Es��ʚn�d�u�۰H��v�q�����qc�4:7�#��ºy� FWM�O���=�� �	��6�d�q.D�-�;��>��I}c�$�_�1��)�R� ���������&R���կ���K>/�Z���9�ض%��r �#�]����E���F�,`W`���(� /l�2N>����k��=�c��<���~�w'S�� J��/��u-R{Ox+Mv�<�o���D����r6�q�5zK� �y<6�mӢ��J�O������>'�?	�,�no�� �E8�*�:6 #�O^5z~lM� VE�J��l5KmI䰷f��/��`�^\�;��@ApI ��HP>\�Kҿ�zw�u=7��VAo��F~k�	]rr@��c�$�%�%����ض���U�<#������<�c;�v��=jy��]I����S��[1[m
��q�rF99��Nv����=��4�AnRQ}k{�M���܏��~T=@�Ov�����%����x�3�=�XS~~�S�6�<?ỿ�Zu��/�I���g͹�I�P�Q��ҹO�+| ���X0 ����W쮔��YZN�����ōqLYi�c�����]��&������Q�w��4� ���Ȯ��3`cq�@��+3ǎ�x�{��X�O����5Z�GKg���R>���d���Hċ�L3�M��^�&I?��ׇ�����n�[�R`���#�
�g�������G;��9JKF�P�h�V���ݩ��G�k�{ӌ;c�yS�[��ZE����ܮ�Q���j+l�}����;V&��Z�s+'��Pk����n���$�yW��U��z���XB9����Qܞ�~8��Mb$�M\��U�kĞ"k�f�[ʷ�Y�iUr{c��� |���ޯww���+�ȾM�L�d$ �p�s�Փ㯊!����x\���Gc	�+�L}y9!}�k뿀?�F��:�A}|"��.ԋ�ݡ���>h�ϿV<�د��Tr�sUK���Τ�N�����x���ކ<_��'�kKȣa���F?k����[�������%%X�H�`��u��3�ʩ$23/A�������O���]>o��� -Gz���x�=���˪�v>h���D�y<�0*v�
�O�Qª͂J�;T�<� �w�=E~�7����RW}�EmJ��Ǆt��x�o�6�Y��O���x9X�
"-�+H����f.ܓ�6j�����I�'�%���߅n����<����^Tc�I�;����"Z�����(ϟ!$t?1�ںk5��V�:�M�����0o�9�d��Ѯ��?��j�n@������Ү���b� �f'Ă\�<�}�*�$��䝣q�C�n,~.iv:��i�+�����$w! �N�ןq\=���=�Ņ�mwn�$�������]
�\���Qv��؉c�FzԞ^�5F�852��p1]NL��H�Tm�Ӄ�H���4�Q�һ3� ��+�@a�9��V�Zz�E��3D:�=��d}:����<MJ;A�o�ՙۤkL6�zE6xdn>���,�$�*��A��� S�5YY����E����bhz��\��<�cΚ�K�䷖b~w�k`0p?�5�� ��������Q����_rc�����S¾*Ӽe�[xGŻ����ePe�n��S�^9�]�e���{��四YM$|��7}H�`�����j��
~�C����zѼ��:�ޟ|L������ܓ�g���g���wg�I.|M��7jm�@�m�69 ��ڙ�MR����,��o�i��}�(e��*{t=+�V�h)����G?�kx�=Q�[(��[3���s���W��e�e7:v�c+G&�?�H*G9 ��5��� <y�[O��M����I�n�V9c-�`�e��\��O�J  �b����^G�4\�� ��?�q��z	�jҮ����5|D�~�^��g�Z�vR�o%��Rn *���sY6�{�xg�z��y>�}:@�\�����<�=k�� f��� /r� �F��"����_�� �u$��h�5jW�9KC���1�w�PWY�R�{�
�\L�\��H�,p� ���k��儩����[�[�$�lu�1� ���,�m��v��#��M�˟ݯ?����t5,H���2�\���\6'��h�c��4F0�ֶ<���w��nǥ�鍧�~�j��q>��j��]�y�L՛�]�Đ<~5N��[U,T��~n���,n���a$h�A�!��㡪�������7E)�:��
���������Eo�ʙ�g�\��GT)]�n��.�O�����z��KZ����̿���;Tך�ʙ�O<u�+�_4� !��T�5�]�J0ۯy%s�1ӯ�C:���5�HӋo����z_�t���D�ܿ�oc�,�����5�富h�n��zM���k*�n-r��FV_0�A��V��߆~-���ˋ�'�H�Ҿ5;bI�<�i�0GC��_dxO��o�]4i�i���Ǚ&8i�^�Z�|�Zs<�9��2v.xSO���-e�ꚋjڄB+��30L#=M~f�7_��uc�`N ��u�{��$�rX�6F�I�k�� �n��kXd���s龫���*����+�4���Y
])��>����J���-�������]�9`Wq���B��%�ç�a�x������?��#����|cᜁ� � ��T����-Ұ0C���]��ξ-�s���S�����C��Q��v�����܏�>@��@��ڻ�GN��.2���y ��ɢ8HS�Y=%#ˮ�:c�O�)�8� ~�d��g���q�zz�2D[>�4�b�K�K.O�@ ��9�)s-55��϶au��d���I� �c��V�t��r>��7����k_A���?�t���*�\)�-#P�WĿ����X�<g�q� md� �i��?���������O�tg� "�sb?�ϖ�}Q7�1�*������J(�$�z�Օ��*�3���?Z��x;T����Kp�6�3O#��}rz��FM�#�R��Y�I����FѪȿ6�º��r��K���4�L2n��0=~fU]C��ƙ�֍-��΀	��ʓ��x���{,3���7�y�҇�zӤV��-��0�D�6p>��=���Q�4��G� v�#�;���ң�lmm��]_}>�|$pH��ℹ��(E�p^*�M[���o}$(���#���ӽ}�o�Bj�e��>��ݬrA"붣z��̬0px�_ G�{T�o�uH�n�m��.#��lIc ��u�r^"���.�a<>Յ���!7��:��}+��Q�F.KS���Ս(Բ?N�>6x��H{�����FY���[ 
���8�9�\��xi:|���eכ����[Fzd�8�k��N���Mgj��"�Չ�fps��{x<Ms��&�ii��u!�I���v����X�#�>�����O�ử�!T��CI+����{�O�����ㆯ�K��\\F��6鶮Ņ����?��ڱ�׉!�/�^|�u߈5� Дu,	��W�����zg�k��j:���~l�|A�G�i%��!R>p2:
�p�M,��8�Z��ʳ��d��w���qi�ݿ��|z�v�YX�:dt!�� �009�}������m�����o�D�9� ��5�P�d�4[���<�NC��춰O
��l���+SO���%�w>��6C$6JW�p���q�2�8��u)�{T0��r�J�=���-Ƶ��ū�joGs ��Y/�
r�Q���ʓR��÷�ͩ�*�[)w���M�rAa_Q�=�o�'�P�ox�A�vSG'f=�pj���I|2��6�o����(�}�?�2}��k/�?/*�fmW�E��s�u˴�<I�_[���s{,��o
��潗�N#��wX�8������O���N�S�N�o->X�#kW�xd��*�	$����X»�'f#�-��?:�U�Ό?�s,/��ׅWͩ��#ԭ�%��^3}:=R� J(,����#������3�^ ��F���"����i8Q�!G�'�w~���F���^-ά"��X�Ɂ�����q߽qZW�Mߌ�{+*�;�pЃ¨$��]p�gR2�M&��J���'���}��󄊺T�'����U����"�#���0ܣ��O_J�����E]WO�h��v�9U��<pFO�T>��Ð�]���m�c�Nra����:���#)a얦u'n�$'�H�ok~X%���oBd>�O�]t��B�L����g���?�/,e��L�������ޅ�y�q�W�����t�.�s�oo��Z��e]*��ɖ�m�8�H��\�c��b�A�)�:�*94	�w�r;�y|���~R�d?�L�!���|���� v���7(皸�X�N�ጳqځ�#nq��ԱJ���1MYW��vMU�W,l[�t���ie.�l�c�N=zr=p�/q���_hԮ�<;��:0ϰ����s�w��?Rqںx���~ݥ��q}'ٞf\쌩��s��x�K��$mu)�#�C�<�T:�����v��<d��[S�����B|H��g�i��c�֧N�}�|���%�/Y$����s��Kៀ���� ��Ʒ��^���Í��8誙�<��\xi��@��a������Ԏ��z�w�t�xEm4���r2"/)�,a���`I����Җ��6�Z*��?���/j�<U
A١ϑa��6���=�y?�l�m���|�JѮ����)��}W��1�+�r��1\ø�l�$��H��RF�#�rN��x���>9�c��Ay����k���Ź\�n�7��j��'�-Ż{�y<Y��;>��4��l\6I<��W�h�-�
�A�^��&����O;?�e�w���p{�^���494I�mWZ��G!&�q��C\��w�|R��8�nU.W���Q"nc��<�sj����P��ԕ�=|I�xK�W��}2�A�>���s��J�v����6��Z���v���L�I#}�ݷs�t�
��ֺn��������J�+9NU���'��V�o�=����Sn�ok��2e�����P�*M[R�Oޮ�2�SL�m���t�p� g�m�ZU�s��V/��X�=oʴ�������'rA�~�Ws7�la���k����|�w��:�1���Կ$"���	%Zs{3Oᖓo�x/E��PM"�f���xܢ��2A#��S���Cᶱ2U1Ơ�B�N=���%��vW���K�����_0��"�1���:s\��%�� f�.ut�k$��Ĉ�H!U��n9�9�z�iڼ�ѥ'�q��>����s�/�+�ҭ�#o�F�-~�Ϯ[Xe(Ypz���V������>tLG�|Em ��Uq_
x�◂������ww��1�񻟿�1���+�~��Y	�Ox㵑��)��\�2L>"r�8�и\��
q��>��?o]:�S� ����E�B�}��ֹ-�� ���t�g�Z�LS�����kO�uH��d�Q���H��?�kQ4/G�?�\[�L�(�	'��@r{`sDx
ݹ��M]׹�v� �Ǌ.'��z�&I�����׏�B��⿌��՞�hn-1��Tl"G��!��	� �>�c4�I����w}�2G��&�ͬ�AKX�rX`�'=�^�����
�wе}Y���\�6�a+c�q���^�ң��p6�(jVU�{��Y'��i� ��&����&�~�=��Ϩ,Com3&�� 4j�����9�[o�{A�����$�CE��~��ڼ����Hb��ancO�����NJ���-�����K�� �l�z�/9��Ҽ�V]GUիz��e�y��g�qhm����(�a�I"�L�����0h�uO	�i�f��Mki"����G	z�+j_�_-�_�x�K�W'��iҮ��ϗ�k����o	��@��þ4�ׅ�4��}��w�-��8ʅp1ң�P�QT�lϙ�L�IB�^�1��OSM��p��בҞ������ա����b�OF(&c���Tnm�9��+�e�I��T�������B�x?|�4|c�����I�?AB�#�Oo��c�E�������v�n^D��9�\�zVG�5��/���ZVS�V�%rb{�W�OZ.=Oz���	t9MK�J���<�3��1��M`������A���?�ax�I�G���F���Z��A-���#�~�����x/��/���wq?�U�nQB���(F=�U�ˣG�ز��Օ�u�3��9������mdHh�_�kֹ�h�_�FI���%�F[ov$ƺo�v�jW�x��c*]J"��'��@����WSZ�}'��gL�#ǖ�T��O_ơ�Z�9�j`@_ƺ����j��(F*#��84��R����+�7�E2�I����JN�2jHcY���bX���*o|@��qu��f+�r�<�3����w�S)�{+��2�y�ogZەu-W�V'����$V�~_Ϊ�����*��b��������6��6�uz�U�!�bA�j���d:����t�U���A�#(a�����ZR��h{�A�3�yR�2ctd� ���r>�pó��+c���ׂ�����:�qU��Yꚼ�z��[�����E�c�a������KO���?Y]���I��8�N�q�mܩ�T�R�y�僔z�|7e:?�W8s�6�C�~���;�\u�x�����ZN�:��ψ"kDU8ڙ�?�A=:��n47��"�xy<��Ofq�qڵ��I��S�J�[㐉��ᏳL��ڲ<��q��Hɼ�I�2x��[�z����,�$�_�Ԉ���WB�q���X� t�y/f�.�^-%��$���Q��#?�L�)&9�:�k�_�_�8khv��^�~�Ҷ�c�>6���qϣ���iW� �֓4���4�7�F�����[>��I��5���x�$������yȪ�\�F�G)���� i\ǥ�Yo?.���=�V��PC�~:6����JˏA{��n��T �?��H����&�eu�Y����]1i���RO+��'=�"����P�,f���Y�;dq���8n(��\W�V�� �ƒ�m����W�ζ�~yU0ͱI ��*[�^������۴�Fh��q�o�����"���ö���,$���J����g�<�;W<p����}K��/dҶ��|^�ܟ㿻�����Qw��I ��<���~��z��Ep�;E�=����/h��*�jO�K�߹�#8��� t�]���(d��O
J���C�ǆ �ϵx� �*t?zQ�Qמ6>�ֿm�^���Z£>h�� Ы�������G������c�h	�� ���x%�ZH��o�*7KmH�ػ�b�!�5k[�"~�f�d����pG�ă������].��6h᭏�'�+y��ڧN�A{]+L�ѯ�-;,���U3���ʼ?ė���RZ^�iӺ�4Ё-��w/ b�t��^�0h�S�r;��<��q��F�>�^� k�|1��DW�f����O_��XJ8�t�{�=xz��>iTI����~מ��;M6���'������:S��*�\H54��?��<9��v�,��� ȵ�0µ�o�^ir��r�8���� ���yG�-(S�ƾv�I��7)Eݞ�<�Ȓ��z��� jo	x�V:n��^�4r&�LY� )�"�Y�x��<��׏5H�J�qH�ʻ|���2v��ٴ}RT���t�mb�2���PA2��+d61�n:������/���[NY�u�f����ޒ\+Ys�X1�:I�8�Y��`�(SVl��08�aRi�v;kM.k����Fl*�3�����>���Z�b�����7p�$P��ѷ�}��'�ÿ�v�0��gcm^��ȆK��-�8��#�wt�
��h��k^$����4ig��|Glp�29'�=+ҏ�5��z}���Gds� Q�^$n�'�V��n#��@�瓑Ӡ�|A�Y�,x�B:N�m��z(��d]�Le����zzb��n����a,$�i�=�跲���9R�,�(��7�{��椎5 �Z��t;��^�#C��m� ��O<֖���\ף�]6�/�$�$�%C�GR~j���J�J2��H���rkN�ݿ��s�h�v���S��8��RZ0m6���X��t�7�I�b�>���r>!?��!� �#��V�w��$]gPm�"�� HoAi����HW��	��-$J�������k�H�!�	%��|����gv����{ﹳ;��KQ��SH� HQ8U����B�)#¦�X ��q��+���������L|#n�+�PS۟����������.��K]U���V��E������Q\
�)V�W�o���-�=�Y�.��h�:�`s��ׄ�;�z�I�>~ht���.�$���nɡ��b�>Lˏ>p�q�Y�z��z't���/��&����~�`t@	)綑��r�(�-r���_A�L$���#���[�t����t�|{�j׾�n�lN��p�4��jӂ	N_��� o���#t��U��*�}P��N�3�tg�%������K;���n0���V$��Dʅ]"�?�]��KLY��rc7�2z*�c�/�J�o���\�d~�G������Ng(eڧK�=q\{��ı�`2�������5������h<O��|�8bDb�F}���:ese��s�2�!��HU�~[��\;�@]fF��_�(���9Y?��[W���_p��FA^>9ۊ�cLG�����"{�5wF�4V��Z{�"i��\ 2=n��
U��/E;�|����
�pӮ)lє�d�V�����؞+yW�Ty��K��[*�7�8}���*�Dҍ�H�.��7-k"�7�Y����/mR�؀n�
N'����R����[ �Q�?��]�wK��j�)�~��?Sj�z��� r���-z�fF A���$ө���4���F͏\�ق=J��5=��o��U0�=
$E�Ꮆq��_�D�i���V�U��y}[F�IX���a~ㄭyj���H2o�X�yD7 V��� ]�3��k4�;`����K�ʞ����`(�����#!���:6~�G�[?ꒊv���������e�J Z�}��d\���x���������50��e��k��ך�HF�|z�'����f�O�V��I�(��d.��bQ�*}} |�Ή�a!ʞ@0�ƿ��9ʋ={>��k E��C�@F
�D�5�7�'���k\�u��6������SS(�#n��Ҽ9*�5�J�w2��̠Rt�<�t�/�Y#�E ����f��W���x,#D�if�d���$R�@���=��^Z.'�X�X#�"���K1��"sO�h�r~����Y�IH�1r�ژ������f���Ʊ;8W�H-���п�'�ST!=�����@F�8�-��>�إ]���(��X��P�9N���?�(+s��wk�q��$�;oe1�T��a:M��آ��ak��ܫA�ؙ�	�r�?y#���00����6����+��#�ε]���ʻOI&i���Υ� NT�rץhȕkur�u6�w��6WrSK����`��7EVoc^�1xP���K���9Yw��i�!�����(<��חy��ˋ�3�n����&���&p��}z�J��zȷ1�>]��'y�C���ӑ7�\aX��?��S���sş�v�+�97:����&��U���I�ᣘ;.?/�#��k�r���3v�,�I���nnY�#�=���+������Vk��*C���7\�}6g���\�7�hx�~=|%�9K��A�PG�19��:����v� B��TtR�7ѻ%�L��zI���ܰ���?�G�Ց7 9�M�c|�jj=e<d���6�.c܊�p�5*����ނ��_� c������tF�7	>JON1�t�Jj{C�Jnc���Ծ6�����$�_q�i�����v�*��ҳ˘�	�QU��������i5+�`���`%�zW�\�Y�< ����a���]r��YP�I�HX
�$�ĝ�U�ˋ�ҺP��)sd[�ߍI�����A�<��Y�R=Vsw�Y펿^���@�[��ԣ������p0��T�`�^���rd�\�`�k�N:���L�$ހ&�D�vr���-(������S�>����`�1^�'D6�`n��ZT�>bukX+��UW;꘥�,��� 7Q�tڷu���$��[i�\�T!~���-3ƻD�U�<����׫��m��z�f��E�M�#9��qn��Ơ-1����ɧ׾�E�m֩�EB����Moy䍑�Ir'EX��j���O�gIC/�W���ʞ��1p���q|�#�g^~��u��&���+� IB�B��Hh�FX���EM������>���4~A^'��rfI�K��>fsE��G���(�W:Y;����&	S��Y�N]Cc@~?�s���H����h缟��[��}^�,���pr
�,%C�I�^�ՔC��ɶ�z��^��x�:�YK��
�D�,��*(���m��H'���P�i�vWYfN�c �d�f���P�|��ɸ��C�V|�Fߣc�N�]9�*$����/��l�����̍��=��������A���w�����7l���W���s�*P=M�f��J��w��d�?Wr�6%GG��v�\��RfD
�>�[�\�M�)\g/hg4�w�ou�R;c���묵,4_����9;�)�T�Y�q�z.�5��y������C^�N��IY��������Z�f�z`E�q��ΧK@���_�ɷc�y��h�h�1�+Bs��8\��9�J�F�K�L^�;��������!wpP����mW�v��l�NUb.e������q��ױ��e�p��f4�d�ޣ����4��B7s��ѯx���0��R4˭���������!�*�5��3��v0��A76��?�޻0Z��^��E��`(��|��d�7�*��p]Q�NM��Y�2`m�-����~�$�N
���ᅥ�Fރ��s��UQ5B��Xԇ*n>a����Ž�̷�sQ��+�̹v<�p��B>��JD��W���U�8�'��w<z�*dg<2卫��������9 Ѕ��0jJ��S<2�������D�4Q��Fq�!;~��>��Zol*
4M���U��[�܆���hL֙H:�M��ѯ������[�����,�9
�I������w�}�m�����3��y�N��[��|Q�|��|I�).��
[�!|
��Vsh�e�MV��aZ������Q� ��'�1.����lh.>�_����Pz,o9_�g��;u����
�۫�o� T�;�{����D�yac�C�`2�_�Θ���_c���W��H�y����N4Y�+޹Wښ�S�@�/�=���f
?��4��Kw��#�C����� -�J��bƀ��B������OY�n���O|.o�{'��,�Ήng�R�h�E��Hs���V��v�������Y��O�(g�^�WO����K�i!~X.�Ʀw{g�dg/�D������~IS(i�iܑ���bw�ޢ�m�8'�IB���
��_���sn��3i���5��غdE3���lo�rS��>�e7]K��_>�A@�Kx_����vy�Hզ�ef�O���m�#k?�[(Hoag?Y�mR�}�̴^�㛝��fV�z� ��\�a�7�9¸=�)�ՠ���Ba�}"5F��Jۭ7�Ľ_�v�'���u�R���RʢF`B��2�v�흱l���<ۧ��
ݯ+ř8@T D �/�KBU��/���D��Ľ}{#�A��'�������p�҇&�Vo|�Ā�uֻ��ǲJ����G���J҄Q뻵6��<��6���,vAw�׾{O�A� *�V�J`�wU����>�?��c���5�`����yXɲ���)�J��5��U�	�&���Aژ��V��o����ţ*���st���bE���1�W���.	ڐKY,���	�ꕶ�R����ⴚ�e*7F��0�#_�,���<��v/�(�
e���.�ݱ�=��v�˴��R��H�()�3K����JU�'� ��Lm�%��!{�X�إ��J��D�5������WI+oWo��v��/S�s����ŦS|��L�w�yuԼ�/(���d%Ll��*$�D�0[��Q;�����q9�eo��������K"c0��@�;�U��7Pe�2e�1�YE�r	��/���kYx3n�$/�4�۳�pN�]y�G�%��|�@��',Ƣ�JzX���(N͸�<6���E�(
(���U|[z>Ng�YŒ�u� �A���ͻ�,P���_�i`4�]��<[	O����s"`2��_.�!��j$ݢq�۷T�5f����y�w[�|Gԟ ���fC|o�+���-�/��"�+y��G��ӌ��:��eK3A<��{O��,��*��Qɨ��6�)��N!.]f�9��$�*a�Zn�)f�ܱ�߯��z���@2�fӐ6��t�n�3H5���w��h6���x�N�%61c䍷����c�����9�Z߼<2a�:����d�3GuI�=��<;�� 
vޞ�b�C]�%V���	H�������Om
HZ}�&Q��X��=^�q�N"�{E6�H��Z����C�S+i�644}�vh>��W�.g�79_7��er^x�"(1
�_�[y�)��ޛӉ7T�;V��C�9�}����;��3>�c�L����~��N�
#�������_!죳n���ku��'S��'7R�$� �m�Bc�(��
�s��A���T�����B���ce��z�>,���:��i[�3k6��7�!�X�����a�$���U|�D�ͨ�Sg  �L��N�K�d��3�X��<���R���Ꝭ&od�H��%	.��)X.���-����.��4�����p���\k�W���+^4�U(1����/�I��%D�; ຄ)Vb�����O��/�A�w�S]��M�δ�^���Dn�5�F+9{z��t��W�sCG� OA�3U��U���tƥͧb]ޢ
g_,�m�Y��D@����u*��}.΁]5�Cz3�'�͖�AF� �����W��7PS`Y{!��bTaa��M�i��o����[�5�l�z߀��U&��������5�<3�I57#¦�!�X�e��S�q���P���_L��ܾ����
�Њ��}�,"t��-!y��]6-�ToȀZ�B��ҝF�-��|�
�a_G��û���lP|ƨ2����S{�b�����ICꍯ.
�w#�)I�C�D�|�
�X�^�9�W~l���~��[���w�.N6�WAp�k���O���h^�]��a�Z��!c�{x��;�I����̷��H�[[��r-f7J�EtS�� uW���1��x,k_��tJ��f���#_�Ǫ,����#�r��Qs׌�Bd�?����}o�r��iKx�����R-��uMq�;���N��*C�L]��8\�ǷތXh�M�c���	�!��{�(��F�"��64������V��a�RךJ|���E/��O˽D��-�����aO̾J�o�|���~�c��c��`��*�G/�ï���/5j����~K?ӯ}��[+���"�>�W*O���»�=���r��3mƮp���(�P}}�ۍ&e���
+R5U2(�=[JzhE 8�����*��f!ݧ:}���-kvt�=��f�Y� �Ŗ��l�6���HD���楨q�9�����鷝�Y����3a5/�'�%��ʡB�\:vdP��e��ò�G�Mh�Q�-�7K����d ��e�O���~�q;��Ǽb���8��Irڴ7@𖺙+6|�P@�<�dS��� �y�����kX@7�����̲��-SxP��d�Hc�[G�N1�f�.,����o��+�O	�c#-5Y6O�)��0���Xp0�{��!��,Z0u,BXdpҍ��>�^|ת��,�!ϛ���?%~䂤�hpK^>�H�@��{��ᙼ+r����1v�D>�4��6��v�����%�V9��0� ���P�t ���n3��\
 *+���Sx�g �_���[�)r_�J�ǣ�����J��g�C<1��z�nL�>�iv�m��g߸�w��6�ZV8���GA�?k�%�����(�SϿ$E�)�[�zsl�+鏭խ}�%\��d-�b��|�$D����ܐta�e_��֛V��]s|:-~Y��(=�=m"��u���_�����ոS�:;�R_����[��8ʷ��>��a��P߭e]u���f�{]{3���;:�.��Ʈ_�1uL��	��?�9�B�E�����t�����dF����މ�q��]��w�z�|s�0i#��8���AR{�o�D@Ib[�Ju+��@ga���m��5�cL%�2���^�2��\:M?[�B�.^�������!0U�s�a��F]��E|Չ��|�5�X�Rx�&�X&p� �(��g}#>�� �*(Y�68�l��������p���$s�B5�/;u𝸭�V㾉��������1U=g\�	'{�=zbHJ�K�u%��%�����b��Bϰ�HnF�no�K�v��j���}���G���Py�WG�9	��s;�#f�{�Ch��sE��tX�?�qx�+�
�]�~C]j�5�D5sb���hc�|��EV׀QjZD}.�Q*�,������t��dW�?���	��xV����5��/>��VRj��`ǂ�7�8�srw��+8���O%EU�}��D@.	𾒴�������p�B1p$E7��';�i��g��x����a'p����*B�A�T9D@dr���[d&*�=�³큧}o�!�ͦ�K���Z*"[V\=��4z޸�e�N�m���H5G�����ʯ�~������v�F�^�ĪGι,5͋,j�^��5v�e���M��`�ԋ�|��L�ʹ)�>P)���7=��Қ:�W��,u��(��� *Cυ�z�)"� �[>�K�6����+;���X_�
)6m�:��������r�,�x�vxm]�,��	��e`#����+Te��B��qSC��V���g�D ��Ğ�mF#-�6(�����c�" ��w�p��ڱ����K�5$��o`B�D@�5=	��[$��p��� �;{2�6h"@�Xh���|��:�5�fz=r��	��x�1-��#c����@S?�x��[�`�ܾx._y*3�#��k_�����RP�>�CQ\�W��e�!��E�Y���'hGD�)��P�`JߖYe�o���{�gy#9u�>H�z'z��P��HvY�Fwtr���@�826�+��|��/��g�'���#��������]�ߤ+ba�.��o�pT}�.����!��w��>��g���X��,1\��������CM�ځ)�எSǾ��׷���eT;!߯&��7�����bt��p�w�~l�|�����1�U)�,���;J�7�@�@�jy �Rm�|���/���27%D�`K�d�=���mS��~��*NX��d���CZ��?��5���/��9�?�n7x���>�"��=^9��X�t�?�^?��I�]��Ůc��	�/<ZY�}[�8�Of;��#�����HZ�����;A��xv"����a%���y�h�e+�d��c��6���!J@-��[�Ԑ֧�<�u�n�[X>�XJ,u������؉��ګ��7v��]8����� 	!ԙ��9�UQ/�D� 5=�����#OP����>f�<�H���Y���l�D]!�u�.��[jV�їqܧ�x�+'��8}\�7$3����!hZ5o���/�c���VY�\2�1o=���o�y�Zإ����8WY��Dn��$)5m��"�1�(@�M�����G���b��fp��$ܔ��n��#v�[�[��i�cȠ��r �>SEͩl[<!ώ�������)��?��$j?`�5��8�D�_P��T�l.�����y ������]PR�3C�����vdz�ֲ��$�Q`D�8��[9�{����	9���A�[�^޲��g0c��3vC'�?�Iő}{
�6"?]d�(��%C�J����
���ʅu�Mb;.���=2��}Z��1�?]�d��N�j�)d��D��В��H��������F���@�)����0d���L��L7/��U���n%	�o������U8�M�9��؁�}zIE*�dM෷��=��Yj1�s4v���{�DٲI
��yj辨�g�/��`Ǯ7��@�L]#G��=D���'"�㩧���|aX�}�ϋ8��aAF�>#�Ii-ט���J����t�����b�	i�ȟ�sN�\W�QI�K�Z.x	��R�΃#���U������&����p.`�=�QcW�7���^�٢��d�X�Ə��{������=R��5WG�:EU�_�a�%�8д]ŋ�����~��KcfD+�-������,��p�@E�U̜5�zF���o�)�W�e��v<�v��<�a��E,s �m�aRr��Ӿ�� ��Az�=��#!._�����k��H�NMFo|��n�\v�r;k���;����Rp��U^��6��~�8�K��5}"@]���A.s]>��2J��©R�k9�D rʷ.G�@�K��V��}1��
L����K~�����	~�Y��W
��W����
5.a�zXӖ����U���z��feEK���gP�OͿSi]���ʖz
�"]��6�(x��_��H7�����͉�ƀ��nf�)xm�dord��)�i�;z��.xb�^9%aRB̄�K�	�%3�T��{^ѯ�Ѩ�D酞Ȟ�h����IGH����e����O��x��f��_�J�N�|W��C3me���[�r3�1����e�9{Ҧ�H��̲Y�(�Z\"�>�;��}��_B�'ĶeL���j���x{Bh�1�j)lt�i�*?hS�.�t�E���/p<��%ϣ��X��+�������z;���Hֹ&R��cG�la�ز����G��k�7���n�8�MY6@u�?Hc������}��z�U�ڎ�;�Q����Wu�Rd���|�]�{�n�.��_�q"�p����{�7�[Y�T��i�7�0��8Y&�6��(9���Z��P3�����)� ��9��`��2l���R� '��~\l�rع�Js]��������S<9�k]�t��j�ʔp2����{1�Y)�G��4ZO�W��ő��u�k�x��Na��)�)�V���s��j'�6�5p0DqT��6x�'�ec1_v ���0����v�H�ޣ�t���1g�DO�i��k��l/�I=�A0�p�-4��_���$���w�Fk�P���䋅Ib-�ܡ&�N}��刀�T�+�@(R>�Df�6����_rMe�=4G�ήK�y��/[GShzF|��h�C>JE��Kǹ�#?���>����,��z����;�|��t����5��όϷRgo���Ӭ��g_<�eM2v��F=r4A�'4lJ��qT���BkËL��B<P٤ٞ>�:׺J��g�u�?W����g%3K%��y�Yu�X�����n�:�x���%|[�8�WʭO.�v��|C6�RG~���H;K3*�s�&~��4��R[n�JK�LO{���r��k���67o���rޯ�>ڱ��Lr��\
߫ԗ~�<$&��TA�'~'/Yi��zt���O��+�;l�KV�R!fȵ�$���y}i��`c�j�����R8zƸ�A)�t���H�a���^�O�vr���3S9W�_���!����J�
1˿���]�y�=��J��+���l2!!�������P���?hv�'�_��&ڤ�낿� dt���q}�>�-�^%�7�/_�!�w���:��4<HR8Zl��X�0	���c�8�Դ3f�d~!��,��S�x�^����Jg��M��P��0y�3���
��2O�6%����Y������}���W߅Dy���
��[��˖�RH�'1�e/��j���Q֊1���s���r��IWʮٜ�Ul��p�{���ZOٳ�[&���-5���E��4���Q��N{��٢�`#��/�K��Py��"�VF?�g:p748ӭ��u���I_����z�M��,[V`)��D]o4٪J'� \Ԙ��˼������Z�ħ��V=H
Xٻ���ڲ]��UG��+�[he&f��e�.��Ȕ�\(��h}���f2�u�Q��x�F�r�����e:5b��*���3�WG+�{m%��D�@v�8��/!<�U�:�P�;L��N]�~�IJ%���x��5�T��o|Wo�y�d�W�#��M*�dDǭ��8,�G6���ڈ&Y�dI����cOFA,�����H]�w1�Mt�|r��_y)c���$]����+M��p5䍊QB��7^�-M��Aȱ�� W#��q''���*$u_���*6��M�R(W�O��F�6���kAc<�ed?Knآ�<��*�h�r�����eY���	����Q��p�#߄�d��
~
�����q؇s�y
j�E���[�?�:�e߼��:zz1�ˌ��hmb}aX���9W��#_�h+[��Y��r����ā�O������X��K`�S���a�gqD��M��:!+h��-����:U?�PT��0��V}�q>�N�j���p�b�o���K͟����Ue���|�f(J���]�Ȳ�U�B���:{b���}�ɵ�Y�v��
`�6Ҽ�5��ʆ_0���:�T]���z�cEr�s>A�ڍf���fTu�)*B�Q���p@�4�� i���n%��g�T�3>`���/-��-�ڐ8�2�����}����X:p�`
���P��*��P�C)��Y�ɐ㵞�P["@W�찔�e1y��y��Ô\��5+�?�ďW��
���e��vn��Sx�?hǅ�H ��W���u-cO巾�e5#�~����5�a��Cj5!�!�!�0�f���OL�Bu��̥�'�(�y�qo���)��M��[S�����9��Ws(j�ոZ�otwQ#���F,5f��<cϬlэ!�	��G�i�'�gNV����<�V�v�`�,���Sw,��+�vgW�po�qH�0�O���k����ڸ�S斑���/x�AS���#߭�B�~xc5e>)�)�y�&�*:I���A�܋{JS�)y��L����rp��m<�i�Ɲ�}�p��ZM��G��pڗ3�OO6���d۟'��V��|��_۬ҪY"kվK�i�m�1%�"��� ��8�&��4��V@6�x݁b���g I�Ju��WÌ�M85�펡��0�×�fbF�/�A�ilyw!Ϛz����*)��xp�?.}���s�d~�!�S�$4K�KӍm���h��*v��!�ϻ��bl疢h���ĀOiqs��y��;tm�i	���I�:�n���@�2�J�Q%�f}���gY�p�ާ�w
�����5�p�{�n�֍�ƿ�19j��d݈0�{C(���v�w��*)gO;]"���׬�߶@4gnW9�Ҕm(����u�>�}ȅ-��N�JH�K%"ȦӔ�vv�^�q^��fi�����[jl��~h��>���?�^�z{s�f�*L�4uE���~ *7��>��{����&y�dw �7Ƞ��u2{�:�-cj}���\�(��h�J`J[UZ�R
�m$\�.aJNN�i��A.���\GߙϤ����_�MGm^����b�o�!�ѕ�ŋ_���x#���,��nC��1A_�=����o��ZH�!�uW��r[���j��[Sj�a�y�Nv���=���0.�����ҸO����� �F�_5ɘ�5��,�NY1��|�( 2k���I��W�zG�f�����͂<-���||��>tR�uO�{��*�:�`֌�;���ɶ��L���3�7*����͡j��)/�vu���W���Zb���"�=���p��?R&Gu���?K6�0��Ւ�#��X^l���[m�J~��iLj/#���]��*���
2��'s����gi�&�ȴ�����˻�h�z�q�q��P(��|1�@9�*�DJ���"ؠt�^�s��3�k'��)���"���Y�!4��|��vHO�"_b�k��ʥ�
���[�n1K���?�ֈ�*�1�9Jpf�1��l�Ǖ�#�cB����g� [�$�i��<��LP�1���$����d$o�(Z�7z��߼1Y�/�h��pG�����\�����ԯ;.��я���m�$�8sd+z�.թ�$P�"Pa��G��憚(�i)�$����J��BEg35���)�tY�^�#T&&��'$�j�ly�����L�}��Ovd�\�Í�rn3n��&z��ߵ�V+0O�l�����C��i����N��>) "4��BT�h)\��ν:6�j[x��~�wNL)ɹ��\�v��k�_}˼�$�5B���Z��敠f#�]Ϗ�g�z��8�%����:���Σ��`������?	"�[��������ݍϫv-O�g`�$�-GNK���V=� r��׬��rLG����S�f��|��f`��ԺC�1�pS�=9���
�^I�}�������*o�K�����b@�������@n������?H@P�䌺z���]���I,�B����T��/��/�M��Nr�+�ŃVY?$��&�<�`T�0�f͸��%�r̈́���#��d1m��j�=���1�m�͛�xE�>�{�@]K6�ʴ�W�����?�,κD�^^�_䦥<��Qk�BU]r��&���@������.fy�S��j��J����/եl�Y��B�/�'�¹��u�}!�#�ck��`.<,����/��;;�9�6i��)���ӬG!�c�Q{w�up��6��%!4���v����]-���Դ���ܷ�&%t����Z,&�7}������|�ʭF	y���i���?��w\e�q����ݦkb�S�W}K�)72՗�[�@$��\�N�gxf��Wb� .#؊9�)�*;���>�n�`$����7�q=YOƖ��*��a���X°�+l��kverQ�g�ؙ�:#0�s~����k6Nt�b(���H�'n6V�ۮ�n{Y�oOI�r�M~x��j�����WM��!�$\G7}:�)����P1^V53컄AH^:�jwup" ����~��G���~��6���ݶ&�"i4+��4�O�$m����q�Fjf�rЌ�{�e���o�����O�r'[7���IQ��13����R� |A&y����H��
��EZ*��q;��k^������7����ʴ�����@:u���邦�]/|�Dn��VF�7z2�]v����GmΘ}�ԙ����3a�"��	���2��Ǡz}*Wl�.4:Я�1�Gv���L��UJ=��ul�&�+��+��=k���F�֏p��T����j|?Tw�40�u�F�;�V�U�a��&��R�ԮcI���r�<�w�z]+Jv�U����W�?�?�MS�Y
iN%�]�IvC���2�\��� ��G#�{�J,����G�UV��l�s�[�Mڙ�q��}�O�L���M���Ʋ��w��.�HS�ل��J�խ>�	J��Pz����>h2Dxbo���K�/������-�V݋��ө��ŗ�uY�6V�o�In�H�H�J�X�����+:�x�5���;V�ӐR�SJ_`Š�Q�<�܂�>�u�Tn�?e�ϸ�Ȉ� S[���>Z`�pU��2��jV|Q^�́j�}�J��	�N�CG�����QD�S�~��}�4r`��e�n$�Td&��]��Б�B�+���?�L�[�K���1s2�?|�����
��9�<)�aT�� λ"��Fs̄�	&A�(5���/�D ��̤���Bh�Ѫzn��y�Zd�W��/����)���Ϻ1���~��ׅ\c�Y����k��JD��o�N�=c��ٲp_���w)���61����uW3��_�rl�~
s�]|^�KÐǥ��*��W�
F]�~��ǩ�@ԟ�&����f�L:U�� ^j?��z@�����"ܡ��F�� �W_��~����.�k�v����l�^:�*A��\���Ҽ5��dC�csm�b!e�]aH$�m���B�O����zZ��r�����wp}����ڤ$�&;��O�ʆ	SI��+<����Q���r$
��ڽ��x�s�M�fՄg@�������Msi�oQdK�]�o��k^�rѼ1��۹\�)~m6,���c�	z��t���R�&�QF�#H�X�P%��B����T�����5%e�e�#��A�%��քBGI_)�������E��rq��\:��	� �� y&�n;ؑ����i���~��5�:�*/&}-���9V���]�8���;��rv!��  ~�Sj�h�`�t|8(�� ���x��t��RΑ���j�58F�m�ﴂ������:��l�1��N_�t�8F�D�ih�
:�������k d���[O����|g��t��w�A�o�jt���ˑD��\�?��	ߘSd�.��ɻ���y�&>�'-���T�����'v
	J��lӅ"��\	Α�L:����>�3���?7���a�.X_+���=֋}d|�~���y��,/S������@��%Н}Ŷ��z�����Ih]	\��SC�M�9^����`�S�k�/�Մ�)�қT,��qb�{-\m��o�Qi����㜶}�\gH�&��BU��	4�D@"�u�e`�M����v/�,#_��9�����[�"��X��a�ӟc��f��=�9p���}~��xjrX|¢uq���đy�
���{<F:נ�hH�X�r���g�yV����Y��I�� ~�Cs��� �]��}0�ü�-�����'�F
~?��������d����`�D�����X�=�3�E �7�����y-80��~Ub�n��nI#�c���^g��e����o,1D���ʶ4���@_)��ǵծ�XTT��h+�p_�����WɊdm��7�OJ	���tM�࣫��� ����,Z���3����$�뮢�O�Rh������X=*���Â���߄�b��(>��R�З�C��P_�����A��~��揲*��{  ��B�,���<�ʪ�}ƮP���Vu\��M���E�1xu1P�`�a��:�C[��,D����$˅�Ų,�N_?�����A�^M��-���D�~��9F�i]]7z(i���N�(�%<It>���C���VP*�Fk���gQW_�1v�R��x�͹"�#�d�������τ��8����4�}�Ed���Lf/���l�4@�i	��}QS����X7����[��A����n�6�<]�]�Ey^O��)�҄�O��&�!�E��=�%�� Po.ձ��`o�dG�<	u2/:*E9h��
���'H@���T��^gY��!�1��t0�Q��V�a��|k�@��4W��M9Rl���N�W���[����M�ۈ��P�wY��8��! �X�˾:�z��s��u���)�~;;{[�(}�//��V"@�J�������D�ɣ�����aD@���B�(�����å�=.	�z���Tv�uw�_g�ֶ��:'jK�+��;��?�Y�}Yd���o��X�lZ��������s�e�	��"���	�$.����n�>��~U���ǽk�xy���{��JB����k�t���9��.γ���z�g���I0l/P�.v��m<�˖�C����3ѝ����ƟG���l�H8�=�/��e��o���,4�ވ%i"��l��y��Q�7�G��k%6�|D�56:orTcU��r�+�nM��e��Rx�1BZ��"W��͜&0	�3${ns5�%��E�\�\��3���0�����"U�g��߲
F����4�f��:�ˆ)#,Y�Zbk��{����5�=����߁cJ.�aίw�	��kv�	s�V���~J5iV	��+]��A�)��:��6/������;)O�RF�z�UO�w���
�!aZ�����7.�^�_�}<��}�=���)1��>a���Z�k����q�Z�tek~��\�:h.-��|Y+��,��Fu�l��ՓJ�µ����.�ҭ��g|V~b�Lc�^���X�Zd����0�T�.2��b����8��F�o�I�4c��b����]��O��+�����m��fgi��=}�i��췻{�?�U�;?�U	�,rbc��w�A��\pȞTM�]u��_%q��u�]�<��! ��V��<f��&.�2d�]$�ys��OH����GzP$�)�����j�gz���z��NZ��	'���\���[�����IX̱��W�YlIƋ2�#:�d-�ܖa���05�E���n��N��O�>�~^���~����r����}{x�*��������j[�s�ȴ%3ZЂ�.�[8�W�T�[�z�9���M�8�����I�\�2
	��L::k��=�[eS�G������:o����Mv��ʛ[��)\�d.6�{�|&Y���a,͚�x �dTs՛�\պ�i�k�%�Dd��� $��Lߵߥfo���_0%��o��]�P9�=�t�AU�<�����]�d �B:��[˥k;1���98���M��S�Q�b�`�����,c����Ѵ�V�CpI��O����0�#=�����8�PJ/B�ډ��r	���	�V�:�[̳���Չ����*��r�]�qR�ܬڼ(K�
Շ~���p��]�B�<���M{��� ���JO}�J%�����{V�ػOڊ��!b���7�y1��#s-��ixxxb�8�����R�bV\���cX�͏cA��EѦ�zs_�Բ�K�;LCV��3���I�Õi��c��J^Bǩ�g~+)/�����0���V����g�I��f��r�?��4�����y��4�D��#;�3��ΰ�1� �[9��Fu�Q�f��I�R�w�j~�iY�k���ye���E����b���s�q>���>�u�Cj�����#=�c_v����PJ!����,�}X�,�o�-�P1~F��:�9He����nz�ҷ{yj���@��LF{`��wdC��z�Pd���x���a�D���!鈱o��[2G����<#�$�#n�S3ǕT!ڃ�:�g�HK��gU��m����-�_����:�K�J��U3�K���}"lH�1���t�x^T"�F��z#���>�S�ƴ�O��aSǉ�Ώ}Ǭ6��:)= ����ؒ�;���m=j��C�oa����Fh�N��K  ��Q�o�z��]���j����t�wk���VN ���9_�=�K٥�&u�����{��u7���}����D���f&6{o|:�"f������>d)C|[���U6O�(�Õٕ�e�Aq`��Gu���j:N����10!�f�i�?e�^q�F�N��Ty�h?����8���v�ZP��O=��h��K������Elw_<gFۥ��tzkU��'0��SFc{߷���,��y���csvA��Zw�8��'���^�֋��sC�J,-R>a�e�Gb?���)#mm��I(bf��NlZ�����\���m�ְ��m�p��[�2�T�&H?DR�G�*�bcۓ����_=QU�N��f4�٤x{`��Ν�J���PƭD���rk�T>�˚zI������GsH�� �ZWH����~8�h�,3K�r����C:\����fd��r>���F��87a���7jhG�1p��E)6i�l��t&�/9ɬ�k��6ᜫӠq��ݚ9M��W���6�PK   �e�X����+  J  /   images/5644ca41-1cf6-484a-bb07-c2f9a6f5b19b.png�WW0 �]-�+D��DM6DKV�Ѣ����Al"�Z���$z����:��V!z�������g�=3w���=�:Z*T��  ����[��E6ٝ�L]�{K@OUco ��� �����|�`>z>k/{ ����x�Z{�xx9��J=  @Sj�r�o3v́�I�L��S�g@`
�\���EG�T<e!�����DʲϘ��|���E-	:3עt�&^7Cx�-��
H%TH��!�U����������C��ח��(���~�|����>��`����e�~�L����E`"#�n�����bng��0�d�w��f��u���R?	X_�B����������`؂v�r��I���ӑ1��ԙ��*3~��_��:a���skZ8��[;��"���� ���p�HZ�������1�d���g/ǚxx���L�	K��%y&�Zt�Q�� PKI�!����O�Z��k�>)�|yX@8ҳ�́ߖ�N��+a�i��?���m�ޢ�[e�O�M�����"si�n�4{f�g��!l�4eqz� 4W �J��(����3=�ͤ�;[AI=�� �Z�G�'�Ci�55���T�eqo�Z�K��T���/���m�p��&�5��(��sց�ѽ��;�:���v��F3��� 氉2��G�;H��1��"�{I6WY�#�JJJZZo����gKJ]����p�Y�*�`��&���i��&�k}pp���F�oʡ�t ���>�x���n�3c�ºk�����Vq�[˛���ai�ɢ�L�7~@�ĩb5�W����`S�O�=�\"�����j��oq[��Z�ޛ��~z�G��/��G��)����Ci�h�k����i{(z��_�zģҕSD�i�����SO���"҉5\�^QY�u��6W-"RoMaJ�`:��󸼝�@�&�GH(��3wkװH<2�wgv�9���>�M(�Ѱܢ�k	u��WKJN>��`�i�꒬����Bfxn'�R��c`P1o�9��T��E̵��h�ޑ�OZO��F~��nL,"�h��UO�����`�}�p�P$v�"%Ʈ�Y7;�>��B��Q�2��'�З��>Q���ߨ�|��>SU &N	�}�C��<&�uDi�ƴ'�5_��i��H��dƱ\�7�[�i�^�6WŊ6G�M*U����o�c|��3��g��4jf4�퀋�Da���B�h�bs�H��Lu���_b}���p��9�ib�h�Hm���I���� ��w~�:�Ǚ��(�Z���iaa��-%�X�0n���4�S�P+ҙ=ߊ����D��BmvI�Mm>���}K��A�U���q���LyKHk&��MjB��}���A�f�)���D}�ü����{����h���xܞJ�tW�&P=�a�kw�m_,#����rׇ�߶<J��V�vg���^���ҵO4 ����l�IGB��L��PS��ڽ�����	�;m�y�}a�.��%\o�jͧ�g�# lF�<���s\RCj�ch.�5O</[ߖR�̔��{o�Zwu��H�UV�E���_�#>��N����1�+��Ġ�E٫�ͺ���vub��Vt���9c�M�j]�򏻏aj�(p$v&�99�r�ئ(��J��Y&躙l��u-�1�}x9��x�=Y��絗�<D���T͢Mxf6���Ȉo�����{�W�������fF��Oʁ�����w�7���C�f�<�{a��ḡ|̴n����*��V̶Q�$��e���YWc8���dO΍��$V� =�z�z��!�Nj��8�H|������~@�����;/4��ʽ}�Btnb��D��WsV�_዁�tPY"ۃ�t�����P��~/�9žcT��bQ�F���n�}kM�F=��(&�����<�{�W���i�1Ӣ3F\QJ�"�i3���%��1�ixjF��aƓ��r�*:H�s�Q�"�@�g�����������$-x��d�۴�D,hO$LDRS{�T����ib�7�G6CK/X���7�ɣ� �)��֚��tWDE��+�9��R�dV\�Ѽ����E���X�;+�[���P�a�Ze�J-s3�~v#sA�;~�sDh	.l�//��ܦ�:�S���Ż��|������ᬹ��FO�����h1 W�f�V��e%����\+C�p��T�8�wʄ1���l�5k�a6�|z��j��������2�zX��:�ϳ9	���P�������@�UlA��0Ԥ����\[j�4�r4�j:UOz����'y)c5�����;�u.S�����t�i��p�*y�0ؾT;bg2015A?�Wj�l��ۢ�$1ye��K�����E�^-����T0���8��� ��p��a
�`h*�Nj`���S�^N���dB�@#�*N�CK����9���R���૕V��v@cy�;�K��z/:�,Xi6S|��궣���M��v]�� &)��\�4���9h����_T����,��u��=�n2�O�R$گ�[?&̽�W���'����>�޸��R��q�ݐsW�t�)���9RqP�`��]�
� }5
B����g	k��g��wf�Hf�1bt��}����8��c�N,���.��)��֩LS ���5���梓EjP�r
|-�������q����F�(���5,�y@� g���Z WMP�;�,8#�]$.%'g�^��!��.�x-z�\��������NQ�{�zAz���Qr�����-wT�1�,T��r��5:}�R��`Ha�ځ_��K��������`��s7}��3���ڑ_�129kzV�0��� ;�#+w7�p�i���L������ xT{�^W(qm���_N@xGY׿�<�F�^�FNz079[WE�D����i5��n����a�Į<�={�ܕ���V�i���ܬ�K��$�GȰ��ץ8IU5�D:9��W�Ռ�,!���%l{)�8Do�P�H�~5(�\@��S�mmu�e�m�ڥs��>+��ڃ	:=s�Cl���Q�X�f	Ǒ�V��a�<Z�5#u&r8▴ ���c����~��?�j����Q�EB���C��C:��h��a��L�І������l�z,.���'1yiV���F?��K��.ϱ����"�lC�&A�{>�v݂���`Ԏ��:���<��Pj(_�q�e�E}��*Sy�ţ��)�E��k�����N>�a��Ȼ�U�Mċys|���_�֕�d�.#pѫ��4d1�&@�h�[�Q�����仚b.��W����M��R�k9�FY=�t�fn<O%����\j�l���t�r+�����Ñ��T�(E�@D�����3jbT��hy��b��A�`j	�\)�v0�	Ăl�r]�_��_�%K��*����d�PS���ſɅ�.��{ӕ�#�X���b�\6��K�g��,id�dQ7�o�|#�p���JN��w��
F�$L���2-x�s��`�
�,"#���ށ��1'Э��x>���
#����-�|a�M��^Zօ�Q����q��>��Ւ����v�Ur ,��[���t���(dN��z*�Vvq��}zR���j�fC�;<he>��4�d�R��f�Jso���|���_����|	.���۷�R1?����#�<=���	�of�d���{�-����k}2`Q�5�����/���q���w���t�B��a�˳� N��%y�{�es!}̰B�crY�	5C���ņ-5+z �!�K��U��9i��hE��������$M:a��Y�UmW���JU������R���)�\�Z�~[O��-#���b���T��\p�������O���h�_�fR��L�����WNs��B����z���{Xc"]���oMe�X-��sī�M�`��E������[���Y�T��0�:������ϟ?�=�
^p�>f��ݚ�4v1>�^���f��"ȴ0��^�f���J�j�M�ZŐS_B�M�/�������c;��[�sCT��#�܆���b���?PK   �h�X��_8
  3
  /   images/57489f55-55cc-4ea4-8258-f1cf3d9c722d.png3
���PNG

   IHDR   d   .   �!�^   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  	�IDATx��\klW>3���?�vR�ql7M���aBih 	�F4��hS���H�

�U���u� ��[�(!IqS�R�j�4&�;i�:[�w׻���|wv���cg/�u�I��uw����{�w�4`H�b濙%�k
�ٟn�N�W�éR6���KCCC�v�����$I��$���|�aM�<p�@ʿ�Al@2vPq�	�L��᠎�jii���2ڲe�,��,��=�}��7�~�o�.>��~��Cs���\AY�)�1::J�XL�c+���b����0E�Q\n`6�?a�Z̜	[w�\��4�
�"���(JB��|>��}\��y���y�j�̝�h��t1 ��������X��rrr�6�������i��̏2�j����ee��UUUTQQ!���A�Xyyy
�(>ȧIp�bA� Q�������w�gQdvk޴��;�oN�G9��9c�ڲ��1��Ջ�x��^E�2�� vݫ���vH*�Y3J#
��Sv�y�F���|
!HT��By,�|�{�1J��i�D��O1ױuT�y|բ��j^ՈcwH�V���RJ��@.i'Iי ��L*H��ͤ�wyh��3�PN�������v�j�**b$}�O���#� 0ہ�����TZZJK�.�lc� �������137~��	�Ht٫ju��+�Q%���3�|��a[Hz�$������Vjnna�֭[iѢE��OD�@�c������������Gn�;�>�Z*�B�QP���u��r¯�����cتjz�p���OИ]�/3_3��_�����0��3�K7!ǝ�xvb4O`η�3��"��V|ְ�y1Q9n�O4M�.]ҷ
�"�"��0�M7� 1�a�$������h�8.o6j�0m�{�<y7P���'�lo&c��Y3���#�1����9,b �:Dzd���drG6� ��O7j��41NG"#�L��Z�4>:zs���H�̤�1�!e�?�>�|��b\�)��{|k����8v�#
`�:��ac.$a1�1Ě����2_$}�`��[�P
b��LwWf!�a	��T.m&� c�
��b��(�1TU�'��nJ#YɎ@" ����I�������@�������7m!�8�m�9XFB�|�]�{�r|����5 �h���T��)�!_���b!L��_YYI۶m�ˮ�>����0�}�k���N�ec>�l�J��'_M�ҫV]UN��������~����w���"d����.^�H�+J� 4���Lit��g�-[�M�����A!�����g�v�|����vwM�I�i��)~�9��(+$g]�k&��+W��,)�U!Z� �"����療��D6`%��� 񋵩��O~�܉?z��G���X ��$)\��˺�|�k �������^��h�����C�O0	h3�w�*w�o�N��p�7�Ap��W>L���p��OJ͗Y_t�|����Q޾ig��o�7=!����?�)z ���ڵ�x �or�Oix��a���YN'k�厰�dG؋��\�ѣGi͚5�v�Zۑ�b	�+ H�����-̳�=��)�03qc�AQT�V�Y# Az{{EZ�������S���&-A���I�:YǬa��|��i��	igS�l�1�Ng��|�t�YA,�Ę���Ux�՜G�W����kMY{� v��g?G��g��lG�$��q��MI&K����l�anX�g\%�*c>�\�<��,�F�)D9����R/��]���q�6� �q���"�W��3_���K��9tn��w�F����6�m�K�u-����`��XS�JЩ���1B�G��������n%w���HԈ����{TRT�R��DR�����yqu�0�G�%^�1k�9���+�]��z��8�̿zK,�~�oJ�EXz_گ���JJ�"�d��@�ŋu�m��wۘv�iqa }|q>�t�q?q��v?�_^�����>0Ԑb���Ⳑ�]�z5����e%Is QN2�3�ļ/Fr�S�_�i YEx�~���2��,c�,� �t�b�!�!������"�z��5Q"&Ǥ��b������ҵ@΀�,��&����s�GI�X�e�(��܈��+A��X�`d���&�dd�/�L{�rB��bx����DVbĳ�R��Ф��7���Q�$eOrр񢧵1,���/��%%%�����l�̉ �P��������K�:���6���Z@�c��.
��=Â��g���O/Y��������]�Q�E�\��46�]̇������6k0'Q�}
�Y�v�+W>��Y�h�U��7���\��� ^��z�ϝ:uj!��9s&�����d�?�`]�ḣ��k��(�ǌ�Qbd����-�Ik�S�l�C��%�KX���Й��%vO�g<���شc�aM�a�}�=�
�7    IEND�B`�PK   �i�X�z��kW S� /   images/65d233e5-7445-4b75-a6a5-2d8c2ad1af28.pngl\	8������)�6S�BDe�ci!{�K��c��j�1C��%{IY���14�>���,������:��L����r?�s?�7s]�Tݹ��v�v�]Rց����u�V��֭ߦ��6�ϫ�m�϶�X��9]��� �
��J=]��׋W]u�\1�]nAF���my�閘��uܘ�A:�)�������~�M6%1hSq�}��z�����H8{�YK�3�;gWF��~�J��L�<<b���FĶ�7����=�90�kD'��޺	�󗾝�|���o�{>��|*�H�3���F�)�> �l������v���9o�����ퟭ�՘ (a�S�@����(Y޼x_�fϚ���h��Y�C��5"0CB\5�[6FGn�`�z'�!���)����!���P&��{=9�Ȅ��p�c֟���|b���Q���2Z���&�쵭c��\.�Z&E�vx%ڳi�V��&�ua�d�x4�p���x���V�$�T2�8���`�I������O;`c��2큈�Hp��G:��m/�s�D��1��ڔ]�Y��&(ƌ2ܔ�"ʿ� _s����g��+�r����[}l����ۮ|{�`���}SsN��Y��^o��ꭖ��[�T�O܊
e�ڽl|��Cm	�	!��t;Vf �Lu�η��1Y?���R�>V��D�1AӬ�LPr��@M�77_!~3�;Ś�㦚��Sm���p䛐~�s�ř���Ե��4�uP��H�/2���˅���L��RC����	CT�ڭ�}�/V���H+ɍ	�Z����Y��q�o�X�%p��-�=Q~�1R�J �y�,	A�	w��o9`��~��,�k7�j?�2�����7��߼�x Y��&�1�j+�Dӟ���%�e{�%؍��_h���3�~�����h�f߂[e��ţ᠝с}|@�ȱ�!�������H���h���aMi8��'͜X��]5�<�ܔ�JUÆ�f�a��//<l�Gb>�P왺�}��W����M�X��9����^O��)�0N���E��a�X��jճ���t�,��q9����� }��"VW�8�ɖ��wn��"�}n�(O�F�	��掤P^��~�Ee�XTu�3��Z�z�s``���u��)Q�\�����"�ڝ�C/qS2=�F���SyZP���
G,YYȳɺ ]�c��lW�k�m�0�q(��B�!���u��R06��K����ГP�l�������w9x��1���1�6)買�ʧ�a�B��v�[83VB[�_�D
��d�z��	�;m`1fWB0ְ�Zޚ|��[�G:�`�L�4�� �/ԍOr�+�4a��l�$� �VvD�V.٩�(8��NX�q�r[F�W𣣣�1:�[a$Bh�vm��wZ^���dاo��˚̌хh���߷oI�l� ��_��*וv.�yqn��Z���7'$_���We��ٿԕ"����c���n�L���{Q�N�sPhg�����ъ���7*Gw��N#���]����w �^��_��|<�a�>!�#���Ѭ��-ܙ&���p��gL�n$�O��tN/c��C6�f �u �,h!�"��c�6ha����V]��-����WK���=1�-T���mE|��֌����v��Љ��Uv݈�؅�.�� �Y���0�r˺��l����@&oIcti1Y��b	!��.qGc-�_3�h5{%��k��3�ru�ϣ/���n'_�7t������7:N�ڭ�[ 	9��(!8V;����Q26�;) �J�7JF��%�6�@��{IFzVق�� z#H*#�*U���3@�1{����Lf��C�%��V�@����	s�}^�C�,`�gřZ�d~/{��S!a�6aq��L�A�=zF�
���r9&o`�� �ֱ���� k��{Y�v��(��9V�7 �"�Eא���u�?�d�m�!c���U���7�Q_����x�p���?����Q�[ܱ5���7,Q"<��+�p癁;O\��[����2A���U!���n����5�bת�B����s޺(2�oK,��T��b�����s^���� ��d���fH��U����8�ZÃY�����W����V\�����U�&�Z�_�����5�=hE.�����N;��TC����;�=�? ̲cs9r�6
-;�J�3dHN�;S���_�������3h8���e
v��%B�HtCV9ޛW�k��ǰY#�%�
�w�6����Yiw�<O\����t����M�ν�7��+P���h����[�1D&��t&�{�A��f�4�+�16�O���tQZ�K+O�ii7[�#�d�3��Oe�f�oT� ��.V	�%��Uh'����=Wq�f�Ww�."
[8&.ʒ9����[�KtQ;8��-O���h�ٞ������-�X�z=�{�d�z,N�$��6�@q��r��R�ws�?�Y��0_)B`­$�8����}�o�no!��1�j���3GG�����s����(���9�/�6ǜA��9��5� g	ģ<�\v�By�:��,Kf���/OKcg��$�9yӴ�cNě���;�7"K��Ey��	���h��H胈Z����n]�����G5|��#�m�-�uQ���O�ޗP�p�UY߅釨�
�=�t�#޽�^��*B�j�-�7��!�R���R��to�\��8�;La6&y��@@�@��*!�U��p�S9��%N ����	-�8/�i�Ä���9�������Y^��	�V�.4g��E�\�0m.��X�W���w�=2����>�_���N ��(
A��RUϑ���	56vw�|��%�a�B,-?Q�'-��DD3�*�G��!�{M�g��g��Y� ��k���x����!N��#�*�1SZ_�ZM__[_��
�5>��M���`1y]T����O�Bz��?d]Kz����"=A/�rL�q8�?��uBǞ�G��,�*�̴�;v�{��bf�U+� c]�N�+p$-Ge���h񹀢d� �h
��]���&�B�(J-n�ĥ���"+.O����a�g��}��Ytt�!�h�s���3�\[!x3&�����&�<[�\�T����{���)N<�����uK��"E��̵�<��$�y��I�w �yԀ���f�z">�yJ'&R;�ptmf����*�:��c#�d�H�8mb�~~ϵV�*������=�666�(~6Pa7�������p(�����h�.�zJ�u����6��D�#�����/��S��8u:$���S�W��wq8ʢ��d=�{���5?����@�3�3����"D�Z׆��<��N(�^üu#��7��u�0�愸�9I��G��Y�+;�G~
7�"5�#{]G����y��+�xBuHJ�A/���J����!�	���"���������޻�7��.�͗�]��9Z�#��a��a�����O2.V�_���� �V�%�H���ח�ii#]�H�N��@����6_	~����y��_TQJ�������9������l�`�3:;����(5�mϟ
keF��
~x`G]]]�jUnjT���J����0�*-}}��T��rWVD��G{�����
,.YZ"���s���y�����S���C�cMX~�ݐ���+�᦯O���)peO!s�,�+��^��$��߶��	�;Ԧ��'|f�Br&����s}5�5��{���-,�����wT�
mVxz��͑p��N�f�8Mc�����"�70(��F��sJ"O,�$ڛ��2!hEl����z0�F���.e� o"��ҧ%%�i�r�3�W"/�a�{Ԣ)�ę����~A&r 쫗ݤ8�������˺2�-Mx�.;��������#&�j�Oo](�M���ɽ&����Sf�s�?䈷�;����W0���=�zy8��
hH���=����
�"�P����x���3ř!Lۥ�Mg�n�5�a���XG�@|rbFA=Trf��Q�+�D"<"n�����5��+�srHh��490H�*-0�HYn�}w4֕�ڧ�������f���Q!'�Y	��9B^��0[<�����m�]�%��%/��U�WxY�bǉ̜��lO��~1��;��h)/�`;L��M�s��hfV,���`���e�����Ak�o�	7Ŏ���c&�
���/&#M� ���"ZvE��L��!��?e��n�t\�<q�8�ۜ�ci�e��vFx��|��1�ʡ�}S.@0�(�<`��b��6+$�;�s�6��Pk��jQ:���e��61��dW���4S�t��f�`%fL|ˏʇ�f�3�ɑ�='E5Z�M۷R!����e`�UՒ��H!�N������uۀ����N��x�� ��U��@y�]xƊ�uk����~�1((��;�5�[#�YF���Ў�|�����������;���и���R����sӌ�׶$'&b�p�8�zJ�҆]���JKkV���3��N��/�4��~t@=X�3�c�xyP�+�bk�X�ױ(w(>��x��_,��q����ZU�;T�D'��,�[ǔ��:��R.<�6F��C�3`��L���C�����z|7�I��s�ʷ_����Q�B_g���u�"vI�ǆ����ol�(�?܋�'쥺{�T���|y.�(�s^v��g�:��A�,����b��h�Dw(��?���C��L�y1� }�@/��S|?ĺO����i��'����C(�IZ�M�W*��Ͳ��mP�+g�^S8-M��m�"�/�G͒v��!�u��*��Q�����$��i;t1g�y	��g����0�0x�E�y�\�"���(�}��6�J��vnE��: 雰�y�u�ף�בPpğm2*R��5���&i2Sc�+�Q%����y�Em`��r�YS��qX���Է�
d9� �?����(++�W-eT����x�� XZZ��EFr�:��BLb/<d[jMKŖ���*,�8���)"��WF��c�a)�8;$S>oB������A��:K�P⭟�C+,v����Hr��%�B:nP���Yx̠k���+S��Oz,?{��l?F��0���FKUg��77Y2��? �ܪ����;�T���Tai݀���� �������zIϲ0�>���g��\��,��_Tg�L<c�g$	H{�ª=@��Z7���we5�&�>561񹈢db���O4
��������K�؈T>4�:--��M��N����VP�^Ɣ]b��e׉_ ��ř�d���a����a~�`�?�~�8a/�"HX��p<�a�%��Be�� X�Z��~�562Z���b�>4�HȰ�M1�c	�����m��^��p��U�'����3%�\c�"B�m{�$��vԘgqq&��r�8~���UNs>�?e0Ն�rs`����?ղdwo�����N�\�T^�j>�e�������~��=�����/��uD�ꯂ�n#�����zOds �� �X,mTD����Dl��2Lj�Dj��T��iY�x���l���E���~��E_��̑T�dt횧#�7��c��x0�����Sü�Y���N%��b�ʣ⷏f�du\��1x<O�Koe��$��_����6?�����eW.Ã�3,��dd\\��?�MH%�Iu����>-敔��t�6�|�'Ӏ)���,vqL$��w6Kʒ�錦љW�� ���)��g)D]`r��"~��[���^⤡�|�'α���|%/˗��GbĢ��=+|�aܿZBO�}��zU��_����eR;�7�c��J|�����/_.�C�f�p`<$\�?����2bθm�ߕ�e��YH`��m�bq�O}lsE_�5�E��cBX�0ؒ��b@���
\%))8���ZJ ��ڃffܲ�%��F�\[' ��[=	]~�C�n|=*���8-5d�-�ie�|�'~�gwP��3�N$flњc�A�*A�j�n��{�O����Ihhx�[�!�������̒�� #yfa�z��K���t5�0��UNY��(T}�1Xm3�RR{D��eWg���T.c�o�n�t
:P� Q��5`:�O�>�A��yj �sDjY���ga�B= B�\?99Y@Ƒ�9JԻI��^�W���p�G�!�?��q��F�G��T+ ��4QЮ³O�`h�J�׮�gٔ��-s���~��@^ǣ��  �=B&K@����m.�e��^��Vr��d���e�̒�οbNn㲰�����Q"�𥳐�LkFF�8������r��Hl�����p<��M:L-��U��������\i�B^�f��J����7����ŵ�������7m'����N�*�1�;��nO�@�&}E��Zt�?K�u��ϧZ�^�F�ߴ�Y�z�e�x�Y���K�4�#'�޶�)�3L}��.v���,i]9f��ȴ]��MO?�)��Q����U@+�z�F�]8��f:�U33������C��Vp�'Nf�����" ��+�4 ��Ox�mX pÓT��gr�R�j�(d74���`;����䕒h�ߢ 	�?�9��9
<K��<E�y�Tb��l/��.B����Ɉ��4�^"X���#�i����Ȱ��"�Յף&O �j,$�♠8�0�����P*�e̶�x�JKC޻�(d?F�4Ѝ�<��fmڞ��f�jeΟV&���$$�>����q� �����@y�ׂEw(4��^������<����I���4��th�[�ŧnU�r����v�rl�Cv�}�Q9/���c��5�vq�AYrH�lzZ�W{E �c������-�z��X������*���b��Ye�G�D]��}~
��t��c��4Sr��:���h@����ZE\:y\L�OE��q�fw�����Y�R����bzT�vr�/<�<:�/�7��
� @�:=R�i�	�D'0�b�+�
�S*!],`d�*}=��͐��w'�ș�׮�>h�b�E >9 4R�(�N=0Z��}���z��y=�+���zZ;��6S�����C2gff�g��Ѽ3��D�*��U%�ޒ�=�A������	�_�a�"O�_�R�C��r�!��O�$��� 
����,,D6�prt�xj5���ȣm��:��z$����ֹ�O���Q��L����G�bۻ� q��Ro�[���߆Wf

*�ӟ�P6Q��=R�ڪ_��D�R���2�G�6��Fu� ����;�DibMC��(��3.+�ҩ]t�cǎ�+}�{��}>�9�lw`P��3�d�϶�ň�[�~���{�h��a<'��u�]����Y+�T���0��Gq�	���xeX����ҵ�'N��\���T�Td���n����BP�i$����Y�ӵ�q����y8�g � U��"�ٶ���?{�%��A���鍖666��~b�3Q� ��Mf&HWb�&h�fʞv3o��rԶu�$�亮Bd���%=����q�1f�����}�EJ��t���¹Ǒ͗j�`CC�|�1(@+=Mt�bm���_)!> e`�v�m��7~����u��ŪIC�A��Jv�E%�Z�[�3�`�o����!���
0�}4d�����=(a�٢S��SFI��S��^�Dt&�f�&BHyo�N�$ߔ:��;88X��Q���0d��(�D9^h���;������x~~�c�VX � !��pt�A�>��ISjZZ	h��C���u��:,��$�a���D:�I�SE�&&���2_o�����q	̫W��4�'0���ȧ�SGȠ�xa�n��ׁB�*��.� .�Ru�e���4������G�uhoT�E���c"$q�+{Ko���(�4w떸�K��I��x���	L/�>PQ};���Cl�J���w����pW\h
�~��x�/Ի��@���,�U�顴�(IG�8�(կ������g�^���
zh!t�Jz�����`Hw0�6�����A�%& \,���8�H��h��L^���iL�]�.<�Vv����ż�<�>�gBs�@O�د'd	l� �3Y0�����u�J؈���L�-=����E��.j����Z��ǣ��&]�Y?���̍���������"e��n@P*�A��a+�@��g��g��
�Wxg8��;��9~66F7g`{G������y|F���b�@��ü�}�hT]�<�%�q�܊C�c[���!��x=�۹�W�>;l+_�o�u�Aj�����{`�9�T��z�XO	}�[��k���쎎�6�á��qa�b+6�bz ����l�.�}����E���x��e�?G��?^��W?X����>ZE�bOT�d�^55�MI�m�����v�&��5��j�b;�������0��0z��i�O���
�����>g�}���,l���!&}%�泇3���z�7z�����>Pw��o!�T�l���*?��cϴP��� ���*�J8���D>֣I�����x
B����N۬�]���X��[=Wq���>�[�h_�2�+�z�H��>p����@;�?�/|>,���;��4���H�|;����X�VVɿ�;9�I(z8٢���M4v߇˜�=-���s��}e�k�a����-�2�Ehkߙ��y>UTTs��	J ��������MoRb�b��܏�$�/jj��V�ɡ$�E
N���<��K^;�����T	{�"�P�M_�GEE���^�G�!���1KMd)�����
]i��6�IW'�����Yp�d�����'hA�h4������8y�L�|=�,�B�G®�c���b���ހ;t�u��Ç{/C��F\�r��c05�1�&+�}�SQds* �q֩����t���oEig.�F�}�P��j�:-�8�]�j} ��S__�q�y�k��\�����3�]Kz4���cZ�������E���� �D���+�59��_�9�,�_�`g`�A�^�4�q��>DL�]F��\8�R���	O�o&f���m���I�f@��2�����a�����0740�=�v���[�f���	!�����s|4H�{���y��:�q���)N�d?P�|�)77L�RoA+��π���\E����z�F3rE+2� =���xv�8�k�{gA���/jK�ƭ5M�ڥ�>��?])����� �Rp�p�:��$���q
�G?�xX�覶������]�����<��#�{ە��w����U�}Pw�cţ��N/Y��F<X�v�������:*g�і���G40�zz Fe۔���4b��\5{L�VQ��4(�N__��� 	$��u��C�/'�n��ID&_Fە^�*��"3����;�y�����CJU���n����P5�_x={N� ���.$7��9n�Z!j�����܄���Hf:���b�]d�Հ��e�G����μc�̵Q��K��`���Y�K�������0���'��n�	]��M�M��ˑ̐�sX��Am�4.K!%F��18"���<�,�عj)�E���13�`̆b�؝��b%X$%@HJܩ�9%Z{KݎTV
X�2!�ݓ�\��B��c�[�[�Ѹ;}���X�f� L��Iu[�5�y��NM(O��h\�Q@��uLQ���
P�?�欄��/#:�K�X�}�Bq�r*�&�N��Fχ�?vw�X.2�x�lx0���_{���ԝ���o`1�O�+fʿ�#�k����!��%��y�f\�r���y��\%_�ڐ�k! �c
C�n���������i(y>Y�?�� P@IIl�,:8��i�FR�C͇�މ��n	x�fa0o�®��3��L��fD`����!�J"���b�%�F�;I������[��r/�9�<����Cӊ_���I�^�Lm�h�7��qn֭�,>�[�E�'Y�V�P�>�?����e	��Vd�����q�	���B4N�wA�A�);���o@-����B7��h�E6P/@��;�s��q���*�/y@x���t�rb�Ū�̟�@Á���E~P��x��M���s+�K�$j'��	$Y��Oo>w�f��?�q�omm��9Ùw^x�y��f;�s<W,x}�j#(�������P{��������K9q�y~o�:kIS׎2~C^���e^~������8�}��%����sU����Y��XW���nzy���/iG!(� ����?_�T������CqV---��3˯��ݼ�U_Z�~�ԃ���x4)e��$��t{8\�7݀���z��F|�U��t�c��O�ə�g5���J;�)�Z~�(�{�*���B��e�F�a�rZoKﭙ�ds֗�/ϘRw���~�>��6s�5�5J\�u�d	2TL���}}��5Ȟ:����VW�8���ɼ�1-?�.�g~P�޶�K�.�
_//92�q���!�,+��NP|��iW�/�2���pnj�Ƞ�,I^�A��N�5%DrʧO���?���7w��SW�����GԚ+����h���Y���^{��e��pb-��Nc\�)V'�̊j��*���;���NAX*��t�/�[=%8 �;��MK�쬍��g������M��N�y�8uܵ;��'�J�;�-~��0�_�e�}��<o<�UDa����70:��>"EБs�X�,C%�}A	�M�v+�͗�I�(���Y�Y��T��A>�=`�:��0�����+>IG䀥^V��*dq����YF᎕E���BJ�4A|�B��3�]6M��`-�<�j��x��=t!0̽�Q�!����$?�a�f��T�Nj���v%$��M-�VVw���D�Su��W�g�/�@Pcrr���
��"����}ư�6�1Z��&i��S�̄�='���~�5v5��HkMá}/+:�����_�q��bRۭ0���m!tD�*�w��{�V/3�êJ^�YRy�&g�"~�nj<�]GRҵX b��Ǒ�V`|�G~u�?��s���2�{^��y����5��i���U�ʳ+�m�@��f�Q'NW,U=�ӎ*N�c��2�0H����zuTG,z���!�"BP;�hf�Ң4S�joo�%�͵;.u�Y�y��LPivLr`���W�G���37&7]�ڵufl���Sa���$�_�Jd�Ȍ���>D�ĒK�[�h��V���v�Μ�-���17r7��;�ſ�?πa���E�,=��^�N��1.1s���S�g֬+�@�����S�:�5w�z~-|���_�+m�ś�(����<��%�-��d��S1Nlz��X¡˽*w��]�e�[b��� ���|���-K /�>c����8/��1����^^�5���M�~�t)��X_�D�����i�ׂjz��g�7s�tR51��Wñ�3;N���Ü�'w� I,���˫UW-o陭r^�-�[���X꟞�B���5�3ҏ�E��~ﯱȐ���*�ݢ�^k�u(|���E�VX����8c��iz�~y&�B�'�(�/}�L�)!>�L4t ��炒�<0��^�7|��mx+X��'�����cE�
Ki{��5K����r�l�����ռ����d,�Mk�����F��R���=&�5��̝n�>#���_B��B|����j.���"��Nȫ�ݚ��Ԭ=ݕ>�rGAlA1��Cj!*�4�k�2df��}��ǘ�>RZ��7��*����	�j��1�����T�-t1�V5ﮞ��r��>r�[��&��m
@����=�"0d� ��jg�����¡��Gy����S�2$U5�lo�����Tҝ�HA5�W�}�"�������t1��qݥO�S��ӮG)�TN7��/7��10�`����l����իJ�gz*��<)�]�o��ȼ�v�����m[p�m�w67�W-=��o�����?��ѴC��ƿL�B�s(���8`^��M����%���A�/��@4Ro=��ߝ�g�����M����^!��;y73콽m�\��
��8+]k�/�}X���ۉb��G�m��e@*gF��x��E$DEޱ�:%����Ö��?�
�,K`��a���:��Lj��{���MW��p��fs�&�Q�m<��3-.��/-h�z��K�ݭ���s�RK�+�����С���.>}��Z�	
W��$��c��P)-�����'��>˒��[G2��AlCm�;���g����2���U�a��B� �*y��M�{�.~��I�i$03��;�?�����Mp�����p%�L�ys��V�#K�a����� ��(5��~	�.��0�-���P��RO�����A�S�,ph%R�{��G8�6��r�A�~��h��vm`sb  U� �q^4j�g=���vϮ߀E!���Lu�Sգ��iY��SA�����ˎ@� 9.�o�d$�	t]~����]@�m����ʯ�n�5^wP-��2E}����S���c]��W ������0p�"�ĉ��ލ���/uL� �,��C�]+�'oԼ�Ez�:�ʢQ�wJ����]W�,ǡ�ns*X���Z��]�vIX k\�NMh�z7�%J5�|��Ӑ%�O�M,.���� ٟ�߃p�����,4����p~�F*^>��^C�P��ϔi5?��G�����@v�ךK#�NU㞺j6˒�-�cj�h���*�ߞZ^��3^*(�1�2Y�ZY0޵��Gk=�扈?.�ݺ"1�x�?�RT���sUO?6����@v���;�~��ʚ���/��֭�!*��5�r{:ְH��Vc��P,9�dK5"��X?
<��?I������ޡO���?�b��N�CC�RDf��e�����@�������\��Rw"�}J��YK��	��\��*f��KŪ���e{7W��[M�NMM��Th+�4-d_��!��>}�ܝ+�`�\��	t��.�(c����X$
_�{��i�ڮD>� �P� W��e�<.��eٝ�R����wD7�3�7�;�'(Bf~��}�gl�u�iA
�\��v@jyF��b��#��y��=�Z�3�j�w�@M�2ҒJ�%�L��?p���=�v%�h�x4����܌<%AJ����}N�O�俻]�2n��	@T<3A�_vb٪�ksg	&k����?p-���")�9��؂��"w�P�R��i	�M>���܇�f�Y:�i�s��A�S��V�u5Ev��^'�ǘ�(�]�5UP�A�x�4JV�x�P�l��}w�[�Ơ�����G-)ZJ?�_5�e]w5jF������0;�ڇ��1�+�z�a������W���D�=������۷��^'��㡖��je�[t�XT�'�ɒQ@�ڝV�RRR�Vw���+�m�u�<�Z�LU$2�t�$����͍����k��Z�V��u9p���-Ч���Js=�����PV�yaV<woP��qepnb�9r�y��
�hq��/��;�g��D�S[��>b~Q��uzX�eG��w�c����ǀ�Ů����GHZ�y���w��/�J��h����c��Zӆ"N.�P$9�ҍ���֩z�y��uF����^�D�M�s0���7����z;�[��E�H���;y�'0=n���e�N�;I��s�XkD	��Pf�6����zc�_�>Lq�5x�]���l��)�5�%���Ji�A6_�^T��X~e"�_�A�ð讪�Ҷ��Kzq5�Ѹz��}�wCG /��Roݐ+,_��]��H%QQ���"�%z�7�82�`�N����J��YNKII�t<�Y�������O��e�*�:�俲��)d<�m����!]x��� -S�s���9!Xr%Lr(�F'�y��r+���������Hϡ�{����^:�Wc�4��!\3�r��K�}�Fz��Pg��$����ч��ʆ�_�̝�J��˹��3a�[�C�;�-HEU1!���49y���{x�E��u*&��BP-R��(��O�J��KccM�δ�߿_T��he��?�>'jK�9�:^i�~&�@A�v�/!)t�����ۈ���F�!&5C�<��.�d\�l�,�K)%U��(�#��3MOtƈ�]5��Cf��1���g�¥�B�]a��˘>6�g���BSw ��W���>���5��a5{�x�f����D�//9��W��:e.�%�y�wTf���+�������_7ȳtAι�*�R,�NܙP��V9���b#��7;��q�M
�����)f�Q�ˈ�E��ϼ:�"���5��Q�rb�'>�K�4V���hm�X1�x���hy�m��AK? ���w�=�m���&k5����K��B���(�Se�Y~���S ���E���bQ�V.���*�"��Q˝����E�H�����O�O������u���]	�{,���._���I������f��E�Sd���6_���!��?!���)�q�%�o���e2)�J��-r�K��B~�����Gi�C�y��z�<V��
^��I�K^/iǉ�]�p	�.�xh�n;$������K����|��_G_�1��^�"�'-�v��3EQ0�v�!�|ya�:� 啘��&Vi����b:�@�_���[=y�G[t&�e��N�}ɢ�]-X[B&��f�u��K3⧫�_hF�Z3U�jn���ǯ49#���G�W�|�+4�R �B}�잵ʬk&����B������Hr��k=Q���1��W��Ay��E�����/ ��rg

�c,�3mZy���5�f�;�[LK�L�.�H�M��U.���B~�d?`i&BQ$yBﲮ_M����@&٣:@V�]��7r>m�!�6"�>�-^��b�����F+����T��d��N}3{#��۠23�,9�������S�xB�s��.��0��5�e�}�3�D}-n�,	�t|��'rW@Ơ�,|p��7�@B��Y��}�w���u�����$m�.S���̭T
�9��~���=O'U�gs��B�ZV�Q���A�k#�A5��;q��3U�ġǬ�nv�1�3�
���Q�{j&Z��~�����σ.�4��j�QT���-�6`�
����N�Oa���������}'�T6>��S#����!"c���\Y���: k���8�I�i	��Cɡ����W|�jز�Z� ��F��ދ��m����?�N1C�?�Uy�K�H.q�~JL�	0vN����k��.?�rQ�݀Z�7Uw^��*�����4ӮT���0�"w|�1��W��4�Q�<�^cc{�$ɿ�5�c��R��!��q�I�¶{)�^a�*>�ⷜ;[�e[�2KB�D�86��bY�,QI����r�9�<A�3�D�\�Y]���d���r�"i��ܞ����P���ѽ���~t���000����8`�l����s<�t���X_~�9� ��,��Sշ]\\��'!�v�m	$?7E@��,�O��'..6ׯ�ksP�<�k쬹Ob�)y��9G�	�~�[Η�"]�wX!�`.�q�z&�+�gvto蝧.%U���wz�K���Mz�z˝�)n5�1��P��Aw謖��S�1��.(`!!���\�|O��>Sm���stR#%��E�',oa}m_<X��jh�=�$1�a5��{���C�����5U7x��~wC�Cx�c�$6���~���l����>���[H��9G)3 �Q�.�Ĵa�^,���#� sz�]��9k�"�KVa�4�'��J�ti��GE���<��a�X�\�
�H��ĈK��w� &�@P���ͬ{�\��l;�-��.~��QhA�R_߃��1"Y.��؃�yjvy�M`����---Z�-��2,�!�˪)i�Ek1�6���lN�Ѥ���K��Td2���By��㫇ʀ5�V���!L�Uy��2899��IcvdLBN�e���( |�,�2̵�í�#��RԻF����zw҃�p�C�|�Ty;�O�8�T&���� �H�1���<�pjBԴ��aYɦ����`���J�K�و�G���[�w�E��RA[� ���ـ��:F1����s���{��s��Ӣ��w���sSw����0��cv����l(����oAl9���������s��h���,�?(�E$���B�7�m�R��W���!����C�T��vөCۊ�
�쵝���>��E�)9�U��Q��7I�G|�c�[Ā�Z��:e!����-5���k�c yA����:m��E:'��PBͿSd�,�f��2[��[��+c��ǵE�t���|�,���]��<p�]��`�j�,4%�6U�U�]=���zA<q3c�����$zt � �=5u�m>1�Y�ŢIB��#���\ș��Hc���բ!c��=0n7�����yY?Uo�ܗ�©pi��1E'�S}A
����F��I&hᆧ�w�4y�N��?� ��@L�<	��b��k*�D2b@�@��K�v�K~5ʨϪ�n+�ȭ)-t��I�
Q.F�?��ԁ�'��S��{�����{8Ĺ6�5�u=�/�eŞI�~p���NV,?�!�*����(��*�@Z���o�=���5~��_M�a@o�O�l�P�/%s�����&1|�9�z���Ʀ����u��v�"�� �u��d#��u��uD���%�^&�X:��O�bǜ��+.��i}�L.�P��\1���`?@�J��!$��k��YI�2�y￠���/7~`Qzh���l��-4�|�O��L�
��8�m� 9�rbפ�?�h�0��4����P�*G)Q��A&[���l���A����G�8���K6^�OwAe�b���'�^a���5�	��Α�`|<��R�e\c�Kwww4y_&� �+�X�sI�}s\���R㷽�33Y�ܽӺ7�8� �m��M�{�<�W�C��q[�ӏ{ �r���o'�?(6&f��!X����Y��.�sC�f ��k�#	��Ho���z��q��H��4avg�N�5������7�BO'�F�?2S��ߖ'���<u��� ���%���2��+�ٟ�r�bD������J�Dd��B>Y����։!��l � ������'2�cVF�,}-`"�=����F�[�O$�%6~|E|v���%g i����@��x�j hh�L7EӴɺ�?455��9�v��/o�}N�Sk��^Ώٱ�������	����RX�U���3Q���Ca�ӹ]�Ļ�>�؜���C��"@y �a~˛�����/ ��i�/�h�,6�>V�S�Ա	��3�ѥȧ�-8�����u�͈�������«{���T��scC0�y���jQ��+K������I���6x��Q?.c�wsž��e��B�� �Ţ��1l�)]%�����'�[:vj��U��c�:���չ������y���D�{��x�	:��zbќ>,@��������%�]��y$̼oC���Q�@s���{�D,GJ��_ю�UZ{������7o��y��ߧ��@�E�n�/���y�~����Q��d<���}��&ngiɫ?���HW�[&2ob��-8/A�FC	9X2k?)��>�����1�x46��������s�/�p�����'� R�m$����/$I�Ѱ�N�	���M|qR�_-'�u2�L%������/�1 �\_�s ������9�\]TTQ�iii���!$$iiP�c萖)%AZZ����v@��n���|���Yo��{��g����qG�G���L�A��������h����������U��Ȗ�C[�~�����Lw	i�i>O9<6Pw��qh�@q�{�ݸ���}#@��3�5��;`x���,,xy"�̿h�`��ź�M�����Z�1 ��W=�����PǺ�<�9"�6F�9]�f���a&
a�o^6�l�&�f����<�8���oj�ނ�y�T=�I�U@�^,����_�)p��PB���]rSC u�G��o�k��Q���/8,-<���e��kN��9ͥ�߆������		,���ee�'�o�Q�DbO�K�N�8U�"�(x'��%	,�y(��	�k����`��A��V��cj�)E���(ތ�t�E�l�z�������ټv-ۄ�)J^t� C�Ϲ6�����x�G���
��2,=G`S�8��#x^��N���i3X�Р�30<c(��r�_�o�ʠs�i�S�-�r?�*h���s���B<�s��گ�fi�֫œ��-{�(�	�r�4@�e#@���:�D���q7�e��9�{�Ü?ȅ�$h��M#��Yl��\��|�����uY����`���7�R<֚������e�cp�΋�ПEL� Ӯ�]���!�/<�%����޼�3���	Qo7�8���`����/��H"@<_w������8��cr�0�<��k���i�y������V�<LqV�����i�O��O��UP����lf���D����F긲��Y^_]�������G���Q%w���ݪT=�3�����j�s��d�?��;P���0��o �pD�KK��(�nRRR����ro�����sj��f�e����y0`�4�V-�c�θ�s�`6[r�s�~U�\�S0Lc�t���M�I���`�V:���$�yG$�-؎��J]����y%��ߏ?�Cޔ�������z�O���|����ޖ$u��Sh�߬���[���=��i�[C̆R!G]�u�5�來��uh��9����߶�i�8%D>���P�~K���r�����u|�~�f�:�e���˵�)��F�32Z�@�����'�1�&��EDDd- kn��3!?��1����:�\��_$�IWfb0�I#e�%��E��cIW�N�!xX� h?���/|����؇Q���d�������5b�R?N�rѧ3���={�+++fs��"�Si.���(:$�qG[����;f�s�� \�ZG�h�앞h�m+Y�A�U�$(����j�w�����Jv��_�@0q��@�����{e澏E��੏ߥA�a銅�e #��c�D"<����7i��,�Q��#0��x�\���ô����C#��,�tu������`S(�X\�(��S@��t
�owt�Y��7+Z8��x+ ��:s:!��ju|ŋ�]���. ] �6a��Ŭ�w�k�<���!~7o��r����3<��O��>J j����\HS�R �&��è��]2e�z>���hF���� -p�*Y�hc+ ��P2V\u��̜C��s��" ;U��lRB�����ّ�0�{���E���;�������������#�7)@�6���M����yͧ��/��};�N=��`:�I�
?8�G���3Z>qU�C�j�x�$�e����D�@�>���#����9�}�,���u-�/DA��k��Z��2/�r�[�b��`�Pfg�-��3�������e,���|�ja�����+�v�H�� 4��Z, ��[�s"����_�>6�ڢ��6�:圣�в'��=���T��v~~WN�_��\H0�
S��M;]����ͷ�`kە�ƧMIM=�-IШ����r�9�fd̑.�{F�Ps����O�ʂ6X�R�c1-���8���d+�OTU$�����;�W�q��y�(Εo�Vˆ�ّ�����J��>!��As��l�������� ���'a�5�9��'�qL_J�a<�$XE�+񱀠�ua��/�����V�sͭAQy0�\v�ӑ��._��liGM׌=�M{�7��8������\z^�� ���@c��hn�6�a��ܯ?ò1]/k���Cw�Z3��Fi_��x��x� #���/�P(��t9�� N� N#~rw)@�
m`]�8��׮�`��А(>rF@����������!��6j3�/?����f6Ld���@�&3�����fYIc�CL���2��
�	(�U8>��-7�����=��J3��k1�l�eE��2�!m�$��:m���.Q�����K>4�D�>�|�NƏ�E�x	=[G��l r�͠���g��to�@�5���|V¥���YE��V����J%s2�%ș0�����b�6d��=_����"|L�|ߘ�B"�N���<���g
�?6�����1�����7o��?۪�4۷!�a�ͦMs� �md�M��;����a�m�	�ww?�5��Z�7U��q?�Ā9/�$��9�5���_]+����+�.*�־n8���&G��[I{I��0D�̓�@Pz�k����]k4�	�~w�ԯ�W��>E�Y��?��y�����g�̠p��`����AN�|KS�fL+3���ȐE��ŪT�f�^��3���M�ZػE!�t�%'"�r���	P!Q�+iѡ��������kP��b�
:7�K�<�r�Wk}�x�"�>Ǜ!�$ }	�cB����e�Aˌ
Y<8���mԾ��gQ �e���@Ҭ��|��!��汽�6��`1�ʢ���c����tO�C_eY_ ���/���UZ���v�r� ��od����!�,BZ�w��_�4Bi]{a�QI����l����V��Ӓ:Ɇ���;[�,B1!8B1�@��
L&i�V�5�~yq�]?��Q�i|� �*�5W�5W�d�=���닧�?6�	�s����-�z��:�Am����>�S��(m�$?`�H�����b4�� ��R�e�@�y.!|O�fLP+�U�^��5?���t����:�	�%�Ķ��א9_�9߫�^3�A	j��+ε���(B���dU ��Gz�	��6[�">����0����Q���5Y+��Ţ�4��,l<En��<���,�2f].�Q:9��5�R�n�u�����GZV�#0M�E�+�(˿7��=�T���OU0΍��,�vu�	FPA� �pw���6��/.����ĩ� �����e/�
b$H�G��"��b��#�,Mܜ�}���:�����W����:��)��C���BB�H�Ж<�l���2�*��f=��.�@%��S}��}���o�Ɵ3�K ���6_7��2)d��e�W�2�	���?�H�9�۰r����o�r��8�(<�ZZZ H���l��Pv�j��l�c8Ŕ��:.L$r�{ �{���n�������Tb]U�Uԕp�dR��d��d8�������g�����X�5���l7G���Oۮ�^����bY�vr�9���#jdr ���0ό�'��vbds�]i��r�)`)�~��g�"��
�H�[�f��.�Ӷ�Ӷ� �j�l�}�C�k�7o[�ڜ������>��ZKꞩ��C\{��uA^��\��;��0N�ȣ���H�@Qx:�Y��!rc�M���b�朆s�bHz�A�C?TL�
y��.j����̊���)���s��f����s�@��8R'ͨJ���@H�� �{$6��Z�o��_�@��?z��Lu���ņ�:�kO�M�����KV<�'!)99�1�UW��\o譱�ɯ�.ɸ�	|�q���k.~*I0���K���,-��+y�\�O(��U���޷o�ހ9�6��%�.5�?��j $V��T�3�333�G�Qc��+�	~	nzA�����ypZ�pNs���d����y���P���"pؐtk�BCC��ۋE#��#��&&&v��"_K�MOp��A�OO�1x��y3��𓷮���u�x{���m@B	U������z/^䲭�	C2&�899�~��N܍�JLL,稡4���$�4;1'4-"��w|s�Di�}�V`����O%�m��_ǝ�JЦ;�s� �M/�"�ܓ��C�꣎�9���=ۿ�a��c��"��"�6�����t�$��h�L�9SGī�;�$F���)�ÎοA�������9c�1&���hS�o�P�>��"�5��*cO��G��B�'Y�<�B�=�j��sr-;c�K/�Rv��7�ɪ�d�ڏw:tj&�s�޽������m�����@�pr�X�� C|��x�C���A�ANs9F��J%�x+��f3�Nj�}Ԩ���1E�H8i�'���>�H��1-��y�$$����f�uϽ^�h��#���Pbq����y4���bc3�=�J�yxi�#�ڄ �i��6����zg�=�E��d�����W0�V<]��ASLz��~ERRqO��3=�r�J^�/էn+;�>�>1B]�o��#�f�b���#"n!�8�z	����hA�������gܓ��՝�Sl���7�9M79�uZǚi���X�S�7(�8�aȻ%ZEk�h���`�/���ʒ�$W��r�c8m�:�	y�r��=�.���}�G�T�+O�9���s�o��X������"�Ⳙ����+�ׄ�Łdb⑱������(B��fS̀���)���'�7�o������o�7��f���ntɕ�6�?<\���׎�~w��Ń� "D���i�zm��$b콘7�%��	��?!X���G��39q!=��9D�R��*��6�&���7��aT=2mԫzĲ��0*����s�J�� )�h�Ua�lz�bQ檅�1y��i�N�;�̔����U�.'�±l�*�&n'M�m�ZU�T�o�%��G��o��~�ج��߁r�g�O��Wh�����I��E�O�D����^|PKL<�n9�����jy�E}�Ӝ��Դ#6æ?	��8�����Z���܈��Ҩ�H�?EWg'����WH1�P�;���X�>��b���H�4}�xv�5�&y��o ��g�S0�C\(�9�zO{TP��р���")�sS'�rw|Í8Rv��Ɲ5�k+%WR����AG��j׵m��bK�~ttD��Z1����f(��e����q���[��*9�	�2	DjFo��8��	d|c�P0d���GY<���c�S;��\�,�j���GO��ku�娍��K��M@���	�#��ǚ���,�q��x��^j��i.�0�{Q�%=���V��J"k�����k�e���ݖ�p�2$Ff�ǝuՃ��Ez��=�;N]Ӎk�I8�$:�#Cj�b�0�T ,��l���𚯽���g9XM���Ǆ|���qky�xrZ���z
���SZI� �zpk�\6�����*���������3�MH�Y:���b��~�q �t�G
�g�sV��b�����bVE3:5��3��q��osoT ��?fSc%~R�����&��?y`�W��KY	��'���`��:�/�ih@�0dƒ*�q@�=��x���Ա�1��7g���C��4r�ȇ������r5x$�f�b��I.�*�qb;��h|�������NR�s�s]�{�%?��i�M4.L���>�][q���늌���u?���AoS�`�}��ڞ�Ƞ쵑�Ww.|p���o>k�80��p%KW��66Tg�����}! �z���_���d��5o0�fг��E��^@�����l簇4|)�G6��\��BZK����D����AxSȒ�n �;1���MT�c_欒��%�����B�Q�����X�V��;x �{�L��\�a��#(J���Yb%��@R�!�u�L�WjA>���.��$��<||�'u�+�����~	�(r2���T�lEV�n�k?;��C�&�����6u��לo
��\k��EG[Y���q���(?����9j!��#������0%f�~:�D��) �bo�>**d��G�
���t�fO�r5��h���q����_�5ߏ̅/�>��U>�4��
&03�y(s	���Ƹ���[��1=�O��^�_���yPݽ{7P% �F���u���ݛ���&����&
#=�L!=񌰬Ť�bsNV����&�>�K�Q�X���q�ˈ� �;o,>^l����%�jf	��F�}����-Z]�������Ӵ�^`�*��4Mo�.�m�uD�B�6����j+�X�*/C-'}�X_g�,�_n�� 1D�@0�Fyq�ؘ�g"��q��u| C(�?�ќa�o��X��1� ��q�tCL�U�����^�b!N��4��de�pV}��>I�(��fDq����7���ap�Av�zɤ0�E�T}ןfC�:b�½R�mI�\�3�A{o���N��wNfpÞ�|�K
&W1����ff�Mlإ�6=�K�|�����Њ��C)�襵���n`�bf�sc��0u��T[�j8C\/���aI�K�I7�Jݹ�B����[ElGw��g(Y�4K��K���h#��/]��/�5�z�z泙�Fnj�i�
�f��A������X��PX��8g/,?]�P�V�0l�xKCd��0y뛛K��ܷ%Tr�Oz.�)��t��Y��O�DOK}�է	)ٖ��b߮R� U� �5����)�=�AE�b0iB���`����	~��Z�G�j�F�ys��j�ʹ#�Ps�u%��]�n��e.����1i^m�25;�h��==�P���R�W_�f�"(���_@�X���O�ZK*,'Q��\t�[�wA�{��-�J��=K
1-7��[��U�83�X�����z\�}r�;Mg�äG�[&옷y�h$�.����NOV� Z�2d:h�z���u�����wX�r�v�j�{���
�IB���XVR�&�.��h�s���ޕ�a7�O�J��u�I
�b�zf���;^�]�zA���~��6Uz����v�vc���[C�=`z11�>>T2�{���lJ&�u������|w��#�a�l�g�q��,T�	L���p�><W%�	s\�]o��'Q�����eɺ��x�����$Z�ӝ��?�9@�>W�V�W�6��2iE��մ�����42<'�yy��������r��KN�
ƭ������z��^�L��.�"�ڵ��:���J	
'��d�S$�}��J	��s����!|�djk5�����T�ٝ� Ȭ�A��6'*��^H�;�̥�����1��܇L����3�qo��8>>	?����{S�"G5�������aītL/������*ʞ�V��@�r�.�@���mZ��ŝ�O��v��7ߓ��88�h`Eȴ'���R8&P������W�#+����.T7�M[E�0�DEp�����G��Y�N���v�"Za!�V���X����#��>$QBw*�av� �)��y�7��s��§��oWgˌ��eG��0���5��'��)��K���<�+��$�RL�H�؞gC�Ƌ�� �:8`� z`b2|�6�8����?4,
���p�ܳZ����|�r�.Y?4��9��;��T�~ػ��l�x�Wb�ԇ'�@��)�PCC5�Ǐi;8���PeՄ�^Z��TVWW_���L"jͨӴ<V�-�2��G����@�g�B\P�~���Ҙa��
l��Pt����y��$V���VzF0�I7joooА���og�Lh+�R�,�^󞪞�Q���J	��u�=@	"�����c//���Q_ᲜBv999c�P��c�����;��##���CM�Ӈ��_;A�,���:XlE�5biF�9&}&+�ǄhQ�]��	QdՌ���j;iE��S��F��[�˪Qtm��PS�%QS��VW�_IEEJ-!�%�B�~Z�]�Pjl���.�c#O��!����X��@���ЮP��8�[���l��(*|e��!\���1��'�>Pm`\VW-���\'�&���-�!���FN���\`�Pĺ*%Ov&�d��p���R$���۷�_��x�ܟӞ/�K��a��啕�5DH7՜_S{ڜY��}=���2�r�̯!�޳=�7{Q��j�l�V��-������l)�,A6�s��=��a0�V4.z:M�c�D 	������j��NJDD��XN�,�����M��\t�푑FA�DFLD�VP6�Uh��������;�h�>Ph|�y�����V3m+��nD�v���Ֆ��Z��ة��Ï��g5�[O��(���	b{>XQ@������yH���t�Aۧ�>��)4!�#_��x�EdA�Px�� �򲲀����X��ZIuM�=�Fޓ��6=�v�����mm����脑]�&s�a�N��<8( ����r���K��K%B��'�v�D3��˯�G.=<�<�p�[��a �g�^�U�s}�����ϯ_� ���/����������>��V����b�������[W�q�C���`��Ai-�(=?eݢyN�,ݖ�4�A��|<m��{����^"H�-=�V�>޲�t� �Ǆ�<������9�(}�#u?�a���)�a2�8�``KƳ�m����9������r';�}cb$��+�.%so����6��g�XX�����0U	榏}s�W�s]D#�aQv�W��{g˯Tn���c��efc&���!=��m kB��1 U�!�<�P�Q뼌U�_��C4��N���б���ۂ��o�o��k�P������4Y��%� ��,9��I�no��}���"�v*p�؉*��{�)��)]��S����ыB�:�P����G�*kj�uc�W5狐g���}L�'sz�XF�Q�@*1��i���{�.j����ۛ���������-�x��}d�y���M�\h��))�}7B�����U�i���x�E4��Ď�gn u�)c{x���6�`6����#���Ij�^q�;�١V�dySS�֖c�'����vI=VF�����qv~��W�2(��s��őZBs�Jkv_{?eQ�2f�=�g��f9�|����|�O��C:I��g2@� �\��>-'�ӢNQm���@?lⲴa$J�=�e�UG�S�$��N�ՠ (��"rPia~͉��$�iRSSuttZAx�s.0�l�?��%]�j����P��,/��,L�.;�>�x����Pe���[T�".�'`�In˝�E�hQGQ���^y�O�@��Ү{t���>�IIIy<X~��*c�A�=�����z��[�ĥ�E*�b�%H����L���}g�ݻ���)y
l.&RA9]a����u;��N��Ha�c��pC�L$ 7
�\+�t��7�
���Z� 
�İ���tB�p`���Tylr{d�}�P��$���O�WG�L���^eCNK�"U��8Ϫ�)D�	���n�?�=7/�UJ^�M�o��q�!Ҧ�mp�)G�k�?��#�mB�#^��	whl�ԗ\����8[�I��Z��oc�s�ޭ(?#5�,�%��w։��:��Y�X����i��<��h�Ҥ[zl g�u�m��*��l�U��_x��Z;�J��`�g�Q��]-y��hQ� �����%lz��.��yr�����d�˳Ci����]KK��:��K	�c{{�����ӛ1��ļIɸ}�4�{LOyJu�s�_�v�N��܈�&1*�{����ŵ�?\���]J�t����k���MvU�.����ۣҖ�[WQ8��|8�� ��:�!s��*B`��\079%����1^�P��
�0j|�RB)���Ŵ`ç�LEl���)��]�,mȰ�܉��΁3�VA�,�'��q*yb_�
�먺�=6��Gw4� ޡ6�k�>�o:/4&�h�R�ۯx˪�HH��3��j�ijj���ε2����i<�{aa�׊�olj��ͳ���)�x�<��BZ򱾓��>)F bґ��<�3C���TVYtO�X�u��,wMMʮ)�O��Q�-SB��uY_���z%�ax�X��dn��fd�ό�X%����4�����h<ӊba�vg�!k�m[�_51e�ñ����iwGZs  �ˀ�b{^�P���,�@n�Ӂg&��c

٧��µJoK��^���*�����·��Z9k�����'���|T��	?=��/|�#>7�`Y///oo>_ �o�^��#�+���H�YOo��C~lQiH����v�2��+1j���ڒ~`q[
!<�޽L���k��x�O�UVVacr����^��6S����R{}u��JC�X�7�w�4�\��!,}�Y/��J�О���&%��"�e��2�2�6f{mb��e��O�J�X����+g·rZ$:n�\4�;�G�k�K
ll�Hѣf���+����7����1P�%�IKK.,,�KM�.���!6&(�6 m���4�ޫ��
G����Z`��2�d�D��d��ɠꤻ�a�*=β���B�dJRuE�<�����v�4�f���R�B1A^M�f	cl0)E�Dk�ǰ��������A<�FwA*�Q!����+�1��hX7�DX:n��ߖ� �%�Us ��<�ܼD~��c�G
�Q`$/���Td�]}��w�!�%N��־xZ7���s�����r�� �a��O
5؁�y��ϊ���[�!��Y�C�޽��֤������~�����p������ϰ8%fߨm�bC�`!�Mr�Q��_t@,�Y�t�!��o�W����j����b�ԭE�|s:��
:��/�H���~���C�]��Ԥ~}M(�-�ua�a�aG��������� Qq��%�	�5�ITc@��ת��|rX��V��%�V��V6{�~��gQ�dhxᡛ�WL*����)��b�w:w����C;�"B}7F��n��Ο�u',t6���� ����ƼM�r�O������:"�S�;�+=��U����z̢�{T}愇^�k�g�;p8��� fww;��lm9,�O��*�ģZ�s�;%���x���t���	�����5���t���w�����G7���j�I_�	:���")�o��~�	���F= ��?��d��C�^}�a�r j�o�r���UO`�7j���.S��u�������̥�����QU��ڍ�Yd�>�-.�����t�ֳ����N-��c�g#�L����(�L��{V��ɍZǟȀ-~�\m�#�Wp�V�v���@JF�S�9<Z8���m���ލ~��g���kv�CC!��R$n�s�@��~$<H�=��g{H�t�)�����gN�߮,tI)�F����f眨���H���x6l�'VZ-! ��>%mB�D�����U˳,$S� �WμΡ@@ɐ�o%��S-�x�-H�wx�)ܽ]�����hl|��S�m�������b�G2+���d}6�ͭ�׊�F�XY�e�Z�oX���;f�8�����xq�:j���bo�thyA/��+u��bn��i����9Vz��?ML��ߋEjz�d/���!T.��j;��n=*B�ݿ?:r����r2�)��,B�NE�s]U����w��#�s�qx����;e��W�E��Ck�<�ct�έ��_2a1f��|�siT9o�0��P�*�h��e��H��9m�YW����VVV���a���Y�xAܺ�m?~0ʏ�[�ŸG4m���O>�D�}`�r58�|��,cWױJ�����D�R��Hyt�M���������3���:j�����T5.�3��.)|ۨ@�����ϟa���3���ʣ���m�<���pV��[F�z�&�5]cx�W��mU o����3�!䘸�(/>^���<)'8Dl��E����	]:G}����C�佅HnS3���w��2P~kkkra��ώ
�b���������c33JJ�@�:k�Q��E�!����������+T�닼�B�_��[�n>a��c\��A���0u~�Y�moG�����_Mےr�\�UWW�/ܧλWS��+Yw�?�v� 6������<��깿�xR�՘G�����#��m%6n����\�+[Ĝ�;K7�S"��ڞ����Bl$ka�#��8�!�kQ�:�@��*�$�Y�oͰ/ ;666i�)W�����~�计y��+�W֛�oƖ��7UmT[Y��^(	���ӡaO�T>�W�
��k}IX����pw3�DŪ�IP��>w��+�Y��4��<�HJ�a[N��fK�g�ߣ�2ݠ�3|P�p)�n�	��3��Үa��`A�|̷>�.tF���n�GV�,5,����.ZS+���"���� }g~�+��hhp���>��&�g9�����ŋܭ��?7�+=�r��p%��ڵ7l9��I�3/����K�����z�"����nwh� @�):��EX��%��Ǐɩ��J���\Vt�q�r���A�xlD�Č�r��Ub����vz����~_ȕ}і2s����)ޮa`Ca�N��.�����LS�u�WY�{܁N45�������L���|u��/N<~��=� �o�*1��0�g�������1J�a�}N�+�����Z��L�\�����<���c�t�9�th�q�E�2��84�#� :����Ʒ��:���bc�LL~��x�͉�ɚ�H�j�*#᭏�M��8�~ό�{���Q:������ַ�]Kd5�H�k��m/E��!�6����TR"�3����Ǔu�"���]�EН?��B,�V���)�����p���afn��k�NNx���<#��ꃄB�G��Hm��
�m�G�Q��0�o�a)��q~�1q�w�*_�f�/;;;Z���˕|�dgss3�(ub��}e0}�m�*?�ۊ�Lf��q����7���C�����2<��Hs$���?h�U7��]p=J[/OW2��zC)q?�q��+���	��{�: �����\]�q�j�^)l��@1"��{���H�JϮa��BT�����"+&��S���[~9그w��k:��o��ю=�{jht���:1���^K�9��6�YD��A��N�e�_��3���J��QJarpq���~�j�<��@�ĵCs�z-Fx�b��KQ��R���ݦ���f���1A�n�BO�κ�Co5j�_��G�F��Q2vm��+F!#*c�����²���uŘ##�~��+�e�H�8���'z��Rq@�O��A{biR�j�(-��w�+mD6��*�����5�հ�rc3���5Åm���=�I���������jh�����5o	=)�����,����S�zAY�Z��Vh��666�"}#�B�����ۗ�N��<!@�@?,92�z�A9A�2�e��w��ú�m�]Xr�0?n��PQ�l��?��& ��!nwӂ�y��JRq	hQ�\���к�7�J}�ț�����N�=��1q9\�l���q��K`Ao�c0��g��3|v����ֶ����_9(�cg*Ǵ|�\�,N�YR���a0rI�S&�%��;��@E¨��-F�����c	IrZ�V�'��ޱ��dK L��̡<J-��3c0��tk<�nc7W���\V[ۻAr��D5U��%�H�t~'40:7
�JX�NF�
Q�����@l�'��YQ�|�za�(��hl2��[��sx{b��1*b{�kk��m��'j�TǢ�F�Vp��Э�p���[����;�##.u�r2#y�6���|0A���󹠕���t���C]�{����GU�r�l�?)#�S�fKT�kh�
-,�2$���~�����Z�K/�%2Ad��y�Y
3@QbH-�Ņ�d×%H�G�:_*@�O������:���]5bw��'u���-QJ̣δ��o���$�l�I�M @�F�F���۔����+��2 6<�]���ſ?Ӊ\�e��[�	����5s+�p���H��Jo��Q�����]�ä�_!>��?���`�%�@�`ra	�8�������Z���3)9�3:�<���,�\Ge��m����-x��<���`��ҼHyAM�3����N�x�^de�]@��	+�NNI�qq������;�(�|V��XvϷ
�-��2������ �����Ez�vPw��PK���3�FZg�Ұ!B�/}F~~J�%X�y�*�*v8�!�b�H)��_΁=m;�.�UV�:_l���X2�~�����VC,���/ ��3y�����Cw��w�{뺊|U��b���]��
l�uu�s>�v?�679�{z��Q٘�zھ}S��r��R�6�cE�v�iO����>,'=�u[S�:,ӌ~~v楡x:G�9#����K��}�?�L��v]����H&T&y������J�E��j?���-�u�tC�t�?����e��vi"nX�Mκ��V1�?�?"T 1���<0�(�q�U��M�ZO��li[6�^�JT�����q�fA���]e�<����#�_�8̤�$ݰ>���h��qnn����b����R�0ȧ�_�04gd�s��D�V�y:��m�с�����Pw�`����?���ܱ�IS`�C-���'V�t�m�onn��y�����F��������
�z�NrU�9ץ�P���Δl�<a%�ێ�g|��������.���(� �n�I#v\i??'��9ꡮU'F���/��Ԝ.(����5\�9ȫ�k��d����#�hq�pϡ�=� ��㈭`�J**^��7-ƭÉJ�H�h�>�#�A�u�EA�9ߜ3��y�2�۾�7��ν��HQ%�L�@�]Z/:��p� FV�cf����]o� ���0Ă-J�cY��}�8�:ګ)XƹAI�+ǹ�eW��{�����u�=,z~U��#}��_S�o߭S̽�ҝO~(�,A�a��u9�~ǫ_y'=���Z�Ft'N��{�����mNH�O��x��>�P��p��]�F{w7�u��A��/2ׇYg�*�u'�ж$aS���{�4�.�>ȵ2uv&5������|��i�3`�#l��k@36-''��OIej���XN�ښ�G��qy8	�i��tli�;����s�p/��_o��kkV����Z��t~�Flcj̜<���v�1������X�єGE�q?�h R�K˧��C�orQ*�[C�R��jHxx�������c�W}6HI����� �A\~*
v�p��Z��xO��������_͎�bz g�1O6�
�b�He4�����A<���\J �ы�Rǌ����y ՗dk!6��C�Hr��m�u�L�0 �_��ƭIBMZ+8��(�B#��65E�Q?�5���5�mJ�u��~�y���o�! ��V����z�[�jB<JK�%��{�n��4!o�9�"��VA�\[s����
,�~��&�{pi��$,7�ϛ\�Ԟ:
N �YW��+F��~���p���87~Yu��^v�3::*-h8�T��%�׆p�	y���2�Ԭ�|��q�VJ��H;ͪ�qZ;��W�-ש-�G㙋�����C:"(����\oLLLo��9%@2���n��h��Rq�"��ߋP� ����9a`����%��?�wl�?$�'�����O������ڡ�;P��F9�b岁�"/,�ʵ \*�
��n��>k�ӫt��\�"�f[â���g�v���3�''B�2t�u�ǆ��=�����Z����[�a��������š_��3$�*BI#M�����瓞?؟�^�\_rl@Cub_szYwy)�١�˕#�O���+?� @ �b�:��s�}��0;x�\��9�4�f#�Uj�4���Z��
�֡6��A���]��OĠ%�}��t����L�C���2U��S�G�:q��_��,Yp��y �����{�i�F��L�/��܉�1h�$J�2h�th�%( ����B*��R�ƞN7���@Ø\n�ڪq�*���FE�)�C/�y"��3�J�Q��N�cl�-~beo�@�ϵ��B�aRj�&�c_B����{�����_�	o))+��85$ JDA�G��5K�Kz�0�~jn���x,���u�q�ş�Ks�����F�$Uz���葹Vͪ)��(�d�9�<2Nr���IvI-�#h ���(�)��_��QFm�u <�����;���|�t
R\��u��U��X���:��r¸<��#����j8l��9��ښ\@�$*�l,Z���:߉�Lׁ-`��~@i�M�����<���\W�Pr`�:{��n9wNpa!���n�4��#�x�"d�-BA-���~��;N���YU�6ŀ���a����q�'��3�#�����"�|/}�iK/u�dJ"�P6��
;JO��l�RA�6���lL�N�/;�n��X��KM\k�!��'��P씦o[��n��X˘@��XJ�S�T�09W󢢢���.�c�NU����m�?�0�닒��Q��q�-�ؿU|]^QA��P-q����:q˴_����5�Hkj�n5^�Y�ت��U��<�¨�í��{������(�ȩ�v����}��=�-�A}l��E���O�Z1�l��p�z����=Mt!p�v�f��=٘�E�B�����Zh-���	�V+�x��`u���'�.���T�<��nw�� ���*�O��t�:Q�E~����=������q3�.�h����{}�U��Ü�Q�A��Q-�[t��a"ژ{P?�B q�X�)`�b�3��>,�N1� �������A�o}�6u��5�\\R��O��;x(�.�:���6�
���~����1XM`�9��<�L�
t��Rt��n����R�z���]��.�uUJ銱���<�ޯT��g8��ed8lBY�ϯӗc��,�	.�@9<8���`'1�c^�X3<�L�HOϢr�S7��M���H3K��˦��F��$Q)҅au�W���f�*��oo� �d���_�0��{�ڑa��v�-��w "ם��t������ro����ʁ�bCH�$G [N���=.���ˁ��ǶZ����Z�4c�݂^ �PQ��}}�?6 �ĝ��v��Z�` �o� �\l)�"�����nnoW�Xxzzf:�U��D��ޯ1)�(9�������( z"d���&�qC���{ѥ��N��P��!#�ƶ^nnn��跱G�t�[�N�WzC�rt��2��v�<�ꅅq�I]�����T�5f�u�/��B�F�v�8��zq~�C�S�����~��O*E�3+��d�:����d���,��JV�&�X9Y!'����3��N�O����ݺ����^���?���y]�4gD$�S�S���;5/��!U�P��_���G�����tx/��Û��撒L��f�3!^Iu����w������1R�we3��L�����t�޸n
���t�ni�MMςQ�s�#S�U�U�
�B���S��7�9���"� ��#1�&&��7g�eˀ�9�iSg[�or�x4�]bΰ��]�\���_A63p���(=h����@~oTK�Ω��K�A����RWQ�ܳAI�5#���}�U?�G��0�ozr%���-%�ס���h�V/i�'�H@4�r�O�n���W�~ax(8��vm�e��{��!�䝝]��r�{�V~��s��!����N�- &��k!/>��(��#i�;Zzx�PSS?�oΘz������ڍ�0Y���(����^oc�,/�c-�$if�M~���9���I��O��)wo4�D�oXC�\<[�Si�ʒ�֣���L���ZYM�t��?�:5�(U��ca�~L�ߊuV���F�%������N�M3���&E���Ӟ�w��M{�����N2.�����ߵ�T�5��{B�r��51�X,��e�>+"{�4hnk[�"��SU[;�����fu$c��}�x�V7��,&tN����}~�jdÉ�[DW��r�,z*?q}Vm����"O�I=������r�E�jz��$��2�|�ϲ�T��p���NxW��e�����{2���z�\P�}�'#g��F�᪥��uJu�"U�7V�p�5��!��m��c���y�s������g�(�g�w���ش��N����̛�j���S��;������D������=��ߩ���'#x�����_}݁۷e�w����߷�rpϮ��G�9�t��,�\Cg9&�a��)�(�:��Pp�#h#�����
�,�TG���H~zT�U�f���c"�^i
JL�q����WyDI��3m�<�H����L	E1w�S��:���/[����kr�k�㔏NZ:������R׈�c�7��<���S��y�������V��n�3G�ܤZqb��㺝z-��?oƺ���T#�[�++ww�A60�
k����R��)�||�=/M�3����ƾK�Z�j��j����m`�ٜ���]H��sG�6b
*-u��Z��s����� �-zއ��-?�w
�>�4y��ڈ�O�C\�r9&�>���Q(��2��ޜZS��F5 �8����Ē�h�ν�>����������M�8(�	}���d�=~��ǿ��&��(Z����Փ���j��j�W�v������J����V�#���KJ ���=�鴏���~6��G��B�:���O��y���H���w%� >l��=�W{�+@K�į3T�ҟ���7=Lޘ3���hrPE��+�3���,(QT!z��f�<l�[�t��aFx��!nr.���\�؅�1;��y�(�B����e+Dh�U�Sn�sƐ,�u,�l64y�gk�g6L��r����ʔZ
H_
�ٹŝ��/P�8S(;���Q\������!M(_��}���Y+�7t234\-�C$R�un�tM��pt�8(z�Y)�ˊ$�`��H5��c���pk�ҫ���]M�%ݷ�KJ��� ���(S����R`[��D�eQUIb�ҍ���֝��-�����:J����ܠ�O��гe���!=]ݠ�%������,�Å���9��FC��:���m��l��`0��YxCo0? 2톎~!%B�i�QK���q./��_x�6+�*4�V�YS��*wGXPJ�QvVf0�6/^�H�Wo��V�m׍W@�Z>����&ϥ�ZH*1��_��6�gA�j����שA�܍�Z�z��LL�~�l �O�T��+l�����GAn�����=d	�����4��gv�r���)]�]��}.d?f��ż�+� z�Z�4ٚ�k8!Q3�t�7Ai ���ŭ! K�.l�26��]�)=�����~���/�
%�����ᎉ�|č�e`H��ݿ�
刿���_��쎴��#���\*ְ�5�4)goo���Orp�[ A��Y:8��$ߑxB���wo�5��z�tbnF|SGG��j����#70��$��I��i�\_���x�v0����i��'K
/KVyMX"�kt��m\��~
����(�:���e���4EΚC�A��L�yp�>��h��Ɏ
��7�!J�I�ַ"~=�.���$�Fyj�8>f�,
o}Q����_��:r�I����x�-96��k$���!�=����g%k�����\�XN{�uC�����Ov]b�p��ۻ���*�n������'�"BB�O�ހ����XPX�lcc�_���,��$nnn>�n=$upt�ep����p'��=�4���xj*c��+�?�����~£r�99U�\��LZ
l4�y��9��v�������*��o'/��0�|4Œ�F�窪Pp1��Y�ć�H���؍����i��������%��v�F�?]�E���hV��X�$�ag�\��p
y���uA��0�n7�	#}�o��.2��z�7g���8���a�ܝ�e�f^2 xc�6�Q41$�2��u�Zyf�zw��%��?�r�@~�6��A�9����A���K�NWRĆ]�LLL���s�J�Z�#77���I���!��������-pj�G�1�(^����((�o`�D�$sA�}�9Ec�e36��E��>�NP��\!��ѩ;�s�m� P�M��vǲ������C�k�� X�F�`�Ι/j��oL8�W�z_=��NI��)h/xq��;7A�ip�SA&���+E ��:�]��f�MA�U5�x�ￖc���A#���l��[oYp�u�U��v�Ks�昲^Եl���<�k�Q��*�����dU�4��F��6`{�p�����z��-�	����IPQ�Z4H��Rn� �J-AZ���4�	�U�A/z9/��!*���.�f��k'f�$V:�w�M~.��3{`{�'*#��_MY_����/�S�2��� ��Q��!r�||<�Y�񦂳���k��|?cu�II��Ys�G�o�b^�j��$�g}�Ζ2Q9L2���҄���E�/���I�!�/��/gəc�#�����W�o)���!w7�7'~�U�LU����!��}t�f>�7��CѺF��}�4�7 #� b��7��b��o>��R9��䝠d� Z����[�5���,e���	e�h΍�P�ߠ�����3�q���a��~�ю<|��	˭��H ���"��䇜����#W��}$�urŷo���Z�q;CAtf'��;�C��N�T}��� ��{1HMI&�O��ё!"<^��2Z�,��~��t[���;���M({�u矷�C*��x�8;WZ'�@9B}�G|�	�6p�����͉�<���%�e:z�4�R�>a��y"I�u�=����VQU�=JpG6�]�6w�i�v�8oP��/�D�����l��͠�Ԡ�:4��E)A��F�Ϻ�q�:	��ng$5�>?�a�f��g�dj��ai:$��ګ����]O��$�o��PGlV���J���ºb����ƿ�P�6���׫jj�z�$�'��Z��L��t�NA��Ҁ�D��l쫑Bubݺ>C�ZǶ���HsO�t,@�Û�ސJ�]rn��q�ҿT��w]�l�H�o�vthq��y��L6� ������7c@�3�	Ys����H��0���&uiF9>��[��]=�`�+;�̾|���O�#[��dāMɀ��!�6���P>eD# !엨��/����o���#���dJЇ��$�/̪�I����Օ��a��(>����p�y#�F�3J���|�����m�ad@r�ZDO�]>��km ���SPP�Z�\�HM~'���D�܈�����5��W)^o�WQ�����eGeD��₸��B��{F�i���_JG��'��w���@�#|0|���3ߊ�;Gѳ�uŜf_%pс�q������P�`�\��TG���n�)=C�5E.�}����WvYοxߴ�XJ���M��=D4�k�e����eb��P��ۤoNMM���*��-��e���N0�q���h�D�@��-��M���h���t��W�C��y�@ڹco����tKp5U�78x�ĝ�6Ո�0I�OP�~�;�g�v��-��绫�7(.�O?{w�o�Q:V���8���n�0o��fhZ���l�ߴP�ֹ��@f�>W?�~���&Whe����3St�H������)"���K#��K��BZ�������L�U>4:�)��;֧�#O�8Y�jz@����Ɔ�8���:Z�!{>�[��/�����l-�E?$BX�
�1V�k��w�k
g	<��,(���,Ҿ��ujjjR5�Qᜁ��{{�� _z;�����#Hy�������/}_E�7"�g|��)��Q��B��������Ǝ�.	�-�'a�0��ܱ�Nf�_�J�*�J(fɫBf�AZiͼ�ͦ����xc����q��`u��[��X�ζ�M��%��FR�,�z't	����-��������A3���+s�+G��Q��M�#�uE�{�&_>mk��o.�3�m�d!#��o{�߿g��WA[�<�UmM:��I�e���s0������ ?�a(������ʊƁWXEN�#�n���6�d��D�3�|�������K��R��9�[s&܌,,�^�{���'B��=yr�+�V?{|�� ����|��n�ЗČ�{ŕ;^g�(�ت�w��!"��;f�j��McY��<^��'{'�
e�6��� �������7.h6��Vn�X;�} ��7�������BY���`�,����z��P	M����s*�F�����Vnኴ�{GE@$��G~��ʳ����!MI�ss;~�(���?y�����uq m�z�j8;^���-&
h��Ð�o��䯍�۩�@�J�ӄ�˚�/����^��_�~��ߎ"9㟪e��T�?�{�;�I@yK��t��CF�BMǭa�O曕��Q3��eƍ���@���Ly*w1����U4t�4��*+&������_�w�ڵ i�h��
�!�bm�v�A�۷�7<�}�Iك~�G�.59�zsQE�����âj*� ����-��?�nL�`���@5Ry��;�EZ�?�2�u��YϿR��7�������g
"l�����ޭ�y�y����y}�T��2e�wyk��L�=����Z~�*�;���6���+�ӎ�w�� (��h���T'�j��C>1qq����9i�gll�c���T�N��+u��)v��p�?SV'�q� �zJ�N���H��[�~L��w�����|���ΨM��'=-	 a�}̗���p8FѤ�d� �G~��I*ŬA�;Y�n;�����-J�y�A;ۿ;>|�H������n{�6��1��5�c�Ӿ<AK�A��h/��:����.[-X�Ŝh�L�hSS�ܤ�=}�S�{	!))���Ь�y�|��sĎ��C��t��E6,@��p2�V����O�^���)�����w�ϝ����HM��U�q�/��0܃��p����g�j�\�|3�c'k���9���O��	���S�B��K<���{��R��:Qέ���޵PJWf�2h�t������~)�_�q�H3[+ʉ/�{�,,,J�~C�/�T�[-X[7VW�˗�omU3фq�o��� �f�4�h�y���7�EPt�xmL��W�>�|,(��#'�g}�)� �羅��\��%4�P�Pͼ+�����`iv��_)~{t��ܥ��z�]Ev�`���MY�}�������}�I���k(�3#D@c��
.&'W��CZ���:ؙ��T^"�9�4{�|�����:S��=����\G|�qG�2jz����!�6֊����$<vvM�ܠ��p�����!�21�^�I�A3A��)2�V����Xη����!�t��#
~�`�ُ�e��}�2q7�b�E{���]��S�Վω/������%�QίE�QK�����/
���|7����N�6ݳ��饌#G����8ۯt���Zn��VH�}aho�O��7m��om�%��S��hMjg�r��Ѭ�����W:I��ލ<�:���@���IWU�E����#-i�s�^x���rF7��2ߏ���#��'���ăa��M�q1��#\�1�>6�"\�xp�D���#�!va,g�i�b�`�mg�U�z;v;�.���.�*}Օ�Έ#��0�����t�{mj�|��Haފ�D������F�F��'���@M�&b��O�u��3�~���hcs�_�q/yV��/k��w��[�k��>�ja�M���h1-t���bSssLi��pJ�Z��'{8Х������zgD��`�ðZ����Μp�$1�M_`��8�h(XQATt	B�Q�]MXb��ܦ�����r�ӯL�0����k�H�z��O���~��k��w� #�C�x�Z�����^��{����P���_�����������r�ƟE����t��=V4O�+�e����N[�n��F�-�Hl���E�jL����#��g�YG+�Q\?�ۊ�7�l�F�@س�������0N�%	0�[�h�,�Կ��w�G�Cr��ozOzv�#w1�m�z�&��~��]����x��ܘR���Q�S���ׁ/��e�ɒb�F�Pe�Qn�!7Ĺϴ�^w��H������^}d���h��l1��{��7"���+[Ϛ�jof��)��h\��zy[���I&eǛ�v�!��/Uu+��݀�d�����D�!��3*5�FՋn2��j�'����l����n?�����M���I.���nכ�w�6ؖwV���w?��r����~#r�Pj�I�5Dt�i��c~C=>Rp��JM�^��/��a\�W7c6�>����"-4��z���j1�|c��@i|ì���w[���U�mA����Ѓ��
�f��/�p=V�a�&�(���q� K����`eV�B�&�U*[�D�!'ߎ�ר�����Ύ���[�I9;5���_l�#$ߛb_g�K'�ښ>m9:����Z��E�tlT^�%wl#��ן�ՆA�dP�N��'��}U:�aJm4 �O&�־Ξ�7�ė��)��>wR���8�49\�U*�V�-��p\3���aG�eA��-5���8i��������^��T<K����4| ���6�c���U\w���2�X�Ʒc�|��;2]�ğQ�F���wo�3��f�g:��D��)�P��=WItH$�I? Ĥ�\��fߥ�O"Eoͪ��z	��G8�K�\eY���[�. �n9��znũ�A�;?{��U�n%��\�_��A��fi)�(t^iY�/���l�<P�%�����B�++�_�z����ꍏ״�T�����_�%�t���o��pnk+�zf��$P�XB�Kgɲ���J=6�8����\���`��ܭ��;0Y=!�����Q�E���6,�J?�O�'��|M۠���T����9s�.��G� vTN��[���,���)x��W�5K<v#�	�^/����o� �^ZI#������.\l�<l��<Q��E�	�@ի�?д�[H�y��ړ�(u?���ޗ��/���Y��v�QX�A0�o�B��4=�_�-�}�~��鹒r�鹋�K�Z��v��ho�b]�%I�Q���(�r���9v�e��	[1�%O�Zt#�{�4��B�f^�'��oCNk���@|5|S�O�dAU�B}�����m�f���_��0%����1����_ט���I�ֈ��v�BQ��]� U��`��_��K�/��T�y������=:IG����y%�
�h<�399�cb�wp�=��wj������@|����:ڞ� )�mjjvU����q����@�efff��(3��Z�@�J˞�)f�;ڢ�΂j��߸U��q�k�W	���r�ڿ��=\��+K����� 66��yFHC�Z������WA�l�1��m����/�0���naE�c:�w|x����+&�Z�+��7{�Nq��+BS&���׹� �9Y�0�I?�|�R%�����P=1��-�[��~��2 �Gn�pw�$X��J��I�ʮ��O�I~i �>\�j�<�a�6a�U�F+Xwv�g��d���_'rꑲ��/�Mwz��; @�[YЕ�����r�ϝg1�?���tr�6�h@'Ѐ��ۚA{c2܍��Z�'��}y;W���/�� 8XI�y�6�^B�Y��x�Y\�p�5�
������컇�t_޿�q�_-��Њ
aA#x٢S�(ғ=��Mf'6�3��-���U�Y�+־���0p�7�w��0�ۓ*�}��ۗuv�G���6n���sL绳x���3 �Y��	��+�>kG@i�k��A�pa�2ئ��PS��O�%��;6�s@����H:|�*ň���i'f;A��^�������V$��������T�𓟪�$ ��*ɨ懐Z��Տ�H)!3�]�\q����
]�O��o=C]�4eo�z���7F�� �Gӑ[�8#�F�G͑М�yu>��#���&��j�x_�oƩS��=Ѥt�b\����$Ü�!����ðں���H���_y$s�E@P�>�`�p�$ ��G�4$�ҥ]/�o�9*�n��Y���/��(�`&(+�%���_��^�!Z�_�wDI�-��!P�h%�Ϻ�Fn�r&�z���X������Y�}~4�F	H�z�Ļ`�$R�\���Qd\A��C�>t�(2������y�^�=I6�Gִ�
\DL�z�C6��P�6 C~��G�S]�c`$�����3�ne�1�-� IMM�A�tρ���D
M�2�	:��l��
ea,,Q��ŉ�:=ԑ��fӷ��U���xQ���k�n-/��	4PK�����#{�\�o�(T�o?����������f���AlYzy����W�
薵@py"e>�Q��+�-ǁ��b�ew,�����=-xZ��ņ]�-���o0z��_I6�~����tX�j
|�o.FJ�C^����_���gB��?�������U�V���a;��`����R�'��-.�A�t�)Z��s��˗3�����A�l"��|
r%K��ԭ�C6]ʋ�&�nL�Bƒi��E���f3wH�C)�?w��bQ� ,Y�W���>X��7��M������jw=����?4WD�
��dxO��M���k�ˍ��M_V���������ysy������#F�#��PfcX��$j4R����a�O`'�<��������JgU�pz�/��@6 �nG�spǹ��[x�R��*@���ܷp{�*��WL���t%��)9�hBZc��0�Ai7�H<Bz�m�zy᧪S!�[��s�@Bis3nxee���񚯒MIR�Ȋ�էH���kM��@�Z�77�5�s������I`��4�D�+pi����uY������@�W;L[fw�������Y��ա�Aӝ�tѿ��`��6b�>��nD|Xk���k�ͤgI�8����� ���S/�oi�Z��v\�x,��K���@�7 E4��F�U:�CG\�PpOo�v�܄[�h��\~���>$�}S-C6��)�yf��3�q��C mႹ���uv:��7�W uo��~/a]��A�W��G����M��@E@̟�9�>į&�r�x�E�8�$1K�t���++�ՙR��ώ�*���]����N��_��i�F��2.��+)�0��k=���}58�Y�����*�Y�.m�Q�U��O�u}��o�l]gR�/(����$c�fB�&'�8��)Y�h,��)�����c;�!�9�����.	����+y��SSC=��5h��x�{4{�g��J'3����7�^��ɔ:1���ُ��*����>҈��M(����e����@qL\�)�@[�h�w�ܯ�+/�O������ؒ���5����p�����~��X���x��2�ߺL�
r��Aruc���X����K��ٙ<��ͣ����d�{���z�I"ef�A:z&�@Uyt$���ns`Z"����ۆ����3����ݍ�lv�ɕN�����,� d}�pC�������&��C�����N׻/.F�C�[�6Z��HS*��kF>��-�����������{M�gl����v�r�R�?55�{��b*���X"�]; ����1���p&:�o719�(����pm��:rȕ_�~2��ۯ�:__��ʴ甑O�ep����Q�#��$���h��U+ ������l�nWQq����H(ğ֚Z�^�j�5;S�f��7����?�+��:{䍺O66��߿�����+0��U��m�����}��s�`i@���X>�N�U�����ѡ�8�0���ƒ�����9��]�z�r��|I�͒�!���q�z���p63w	�`� �����9���Q�����F��:���<I3%tyrk�f�&��I?��<�
��_ؽ/����%}"�Z<�A�E�^��N#�h���ޘ��Ml���{�++/���OՅT�_Y�kH��(�(=dF<��Z�x�g������f�y�۸��M��WB���e-?��d`a��u���0�A�����$=��3j�_�_y���`�PŤ7����|C�k\w�����ǈ8p1��n�rW����C�CKbw�i�5D��V�|B�v%�ges����6{���[V����=��+��(7�pӅ�Kt�� �g؉ع�����#*-��U��c��k���|����[�d�[�IO��-�?��f'ʯ�����������J�3�#+����Ϡb��0��ǆ
��t�h1̮��'_�KP�Kh�/$W�]C�Y�O�'�+��$ӑtË���'NlLL�X�Zi��P�a b������G���>��7r6���]��u3��o,HWe��Sn�_]�2Vl%�@�~A�3��w�"3qv22�	���y/���ex}�֣L�hL��e��L $��Kc�u{�F���23U���@��)�K�鞪���P�G|xƃ�{}o:�v���)�X!W�6~��a�����l�R��_�L����3K&��ZkF�݁<�F��0(�K����������H��&�}#r�}Y�k�5��Չoa�0@�5.&�u����
w�
�OPs&&&����|Yn&X�;��
%��G#x�c��4�	�bz{{e�=�YJw����/A�Z����������F ��B�0I�˃���g_�"�y\�h��L��WB�X��b��K�DB��ȕ��7��~[-Xk����K�h�9�&�V�(٭6O8$�n\�ǿ��9��eR@䭧�L��������i�0��zǴ����D* ��K�I0e_}��	��ʁ�A�z&�����)��q�Yy,�J$~m�phO<�ĵ&�W��Uc����Հ����x=��{ʵ�>$b &���7V�#�l63-1%i*���� ޫ����n�@�T}�E�w�!C����zo�6�q�J�� ���S�8�`��7M����.؏��L�O$�/���3�]H¿l��F�No��A�Tƹ�����d�W|�/17Ͽ�Q�|=�����X�r�W0�`%%]s�V�S=�nQC���[�ã�[�k4V�u�6���w��	[GՋ���ä֚������Km����~�S�8t�453��H���������93����k��7�76�~��fZ������cn(�WW�Ժ��,B����ԷWݷ��������<�F���;#���q�pY[�f����g�N��������;���6��o-=�	$H��Bl��g||�r1A&���S`	�	��d׮�m�����.cs� �����&���+�^%��
Y�Ɖq�\�&��0Ծu�NglT=C���T�C�Z����S(@�g..?��ֿ<�����]�$ВL�¯���sQE��oZZZ����J�S��B8Eܵ���NM&�\Aw��I�w��yȖ��Ү���	���W�"�߬��L�H�����گ��r'�"���;V6;x�.A��J��倲I�z��!,ֆy�T��Zc�b���\�ߪ�R�+Ap���χ��S�����K�֘^��l�L�F		І��bP��n��>G�q�����{�æ���F��"w��g��o�]���#[�m��C��/|a>�a��+����\H�-�i�	�u�O����iHZ*�*� Ɨg�k��?�!�6g��"�"�����:e��'�����)rY�/��f�:�E��{������~������}����B:�S��y�~�+�,�2 ��2�Y��"��ӵ�ySl�|�-\z�����,I�V�0XV}x�')��˪p����,� o9@�y}jf������8&��u�+��ԧۗ�Ī/�mO��{*�u/�D��Z��2�G۞|��-�0��CF��!��%'?�u!#����+m��eg�65P�_U�F˗��������Q�Vc�P����5鑰6VII`b����XYY_��n��f2��ň��#�S)6�pe��,����EX��YA�f�2�0p5�'""�"P#���iN1��2�b6�e> �E��H�@"�	��)���d�K�/qw�>-�~��Ȟ�ma﨩u���^^p�}/��=�$�Ϙ/������5�b�60� ��l��ek?'_�fQ��G-��= 5��PuY�7V�?�m��͏ؒ`��EdM	�x����Dw�t� >�t�T{��$�E���;K,�>�-x���B�p=K{�����C{?0�8j�����6/q�����g�P�����H��?5ݗ8�)��~�2�,�=k#��q;�a���K�Pr��|Z������yf���7��c!�^��3�ךM����os;��zv�н�i#?���m?�A�'��������W�"P�j���%%�l2n�ۇ��u��;��@0J�k���$��E��op���@-�d�t�pk��~`�����/1<����^c���⠞��q@E+�Q���+�1Ar�����y7��O*��c6=�JB"�l��Y�S�@-H� ��!�[�P���w���z��(��Y�v������.��Si\�K�̅�8U�`bӌ�@��=v����yZ�~�ݰp��|}A/gk(###�v�蠲Յ��&��1~:*��LKr	�u�k�
*���`f\���y����\�͕b�X�ꃯ�bb��A���N΄c}�c7,U<H�2C�D},�u ��!���b�?���I֭�1��|n��*V
��a�k�]�Y�2�6q��A�/��@0J��
�������u�Fpr���`�K�T8�H��˘v� � m�q
���"!���5���8n��{ԯvY�?Rz��L�g�s�#J�Vo)>���r�]V�=�b���/<d{�YL�7I�W�7���Hā���A�b�����9n�žB 2�&H|���D��cC����)-�]�jJ��׺���X�W\�v�~ΰ�KȩyC2���6?��tK��V��%����M����1qq�����1��&z�o(�}Kd����/���ڣ*�:B���g�6��@`zu- ZP�H���k�\�z�<ގ�f�CN�z��Ý��ʕ��*��~#O��<^�9J���6`��c�N>}[�0�*��*����Ҹz~�o���o��YT��q�kiӶeVb/e>����@�v�� �u�1H��rD����[�3���h���߿PK�^�ZȌd�5󩱤5��V�f8&�=H�,!<�ɞ��;w3k���B��؆��`zh�;G�g�$�ذ�����D����I��������Nn�|�3i?������ʩ�R�Ɗ�:Y�|�{��K�s �@g�#{6i��{��f���[���^�������
���ȇS\������,@GQ1֤�K�������2���Hj�i���{S�/}2�h�YT����q�'��}�V@��g�ѯj5�5a��e"U�����%�D@mg!��%��^n�M{�D'�#	���Y���T�'կj��a����"sF�c:����"z����f�,%%���)�7�b��U2Cdbs���K��l���f�c��&�B�Ly�<9��F8Qz��m�oߊ2»~���>��I�6�*J�f�ky���p4Q,�h=q�!�r���&�(.��b\���yh ;"7�L��wZ�ڤ��5�E���٠��N��myu��q����[&�ZJ�Z�Wc�ZT ��cp�X�SӋ�l��pJ�Z�sVz:����o����}	Wց�QOI(*���UV��_�i-���n��x�nV��i�����ɤ�5322���:E]S�(�K��D[b��)���%xM��U0�do�lCX��|gdwOSm�O���U=�u�oy��]���/.�B���r�����ϵK�������F�du��Ӝ2�7�l�X�U�"��X�����o�������'���J�dK�ފ�YXG�-��ک�k&q���ԴO�p�bk��	�i�ڄ=�#�����������~V´H>��������69���x���ʠK��]��ec$6���wC?=��Ez9,���uvͬ�*��Q��NoJ�͌G�����
蒲o��U�q�O��f6��zH��3��H�.tr�ʅ�ޏ�Ԅ����٦���Q g�w�<�}fcc3��!��";i$�[��RNS�"���������yx�s<�a��1�0�rx��!��X����GvjcP,Hɰ����:�:�n�B�f��2���`��(�	Cn�
��.n ����[b��x7$B� ~��G��B]M�u��kȳ�\p�f��x����i�1f��D�:�u����oV�]�u����ݵ�{\�����y�J��>LUF����U:ؽ�u��2�ZZ9�����ks�����{M��Y�ҙ�_��)��r�	j7mC���4$��:��zOW[����7�܄C΍�"�8ȯ_o!�a�]ⶣ���!Y?�\t�۠A�"ԃ=ơ�>�+Q�>�+T�&��="��9W`�Y���*�6���nj��q�l�Ծt����-���/����&!w	I`L�A�E�iQ�6�o���x<����$!!����p��6JL��gK��3��H������B&Hk7.J������N+�PE��K��?~�0��ѭ�x\�=}҅������S����i3��]מ''�7��3����ӭ��ٳ��-�LC��X4]��GZ׮_��˓5��~��(&�f�!��tX�U�ș��[�!���<��>�f_�v �u�z�z���������lI�,z��KV��3�x֦�$���f��_����:e��	seW��&�,5����

No=ͦq]vD_�V�i���2#���A�Ѳ��M`	���7sҼI���֔�Q�$�g���K����ӍD{YYY���z��i�#>d��f=o���M�r���Q(&c�Kex3���h����|�5rs�g��o��_�]��f��ڮ���k�i�d'�Lq���Ϩ�o�,��p��۞���H�/]����5��3�3���h��p1{	8��	��v�V>>��:<�J{�y���a&�LЁ2�{e�����,>���|�{�<s)c���A��Hu���U���:�����tUYK�ߟ�U�E4�f�v+Og�t<C�Ҕ��Ѵ�!�~�Oo��Z`���x��<�}�2�����妊�ñ}�Y\f&ky`�BҴ��Q��dE����im-fdD��ib"�z�߾,���1%�&s�B�c�p��W\�1��#%G�c�R���B=Y��?���z �8�����Fi�)oiɣ�d�GR\���öp�����p�RǓ�p:���|�ȸ^F��n4�[�����.����T����^%���955�^�(@�1�ۻ�j�w�Nd���1ռ�9&�*K���4.q�/JIr�C+�ݴS?|�"�\����͆/Kq��{�q����.>4�
o\.�)�����]���~uӶJP�g�q�-�&i/�X��F�%A���=�ா����B�4� �6t&��䓞3�uP��u{)�3�>��so?���@C�O\i�s�Fd]Պ'�7��	S�B���B099ycվ���ߎoو�rT��>P:�TQQ��~uMW8exz���56&��n���3�[�φ�8����V���/:e�7	Q���;������́���㑴�3���y�,��@���Dih���i��+D�蘾3��yG��2]96��y��VB�6gQ�R0wu��G�Hb�b�N��w�Y��ل���Yz��o
�Iժd"^���oB��,��%�WיB��.j��� l�k^X���J�8#�O3�BMN�t\���Ƿ��}jf���8`������輟1��y���y;y�	�Xݐ���u��ϧρ�6�?��trQ4��a� � ��Y|������&	c�� GB�s����	�����*����%���۵!"$⭖�Ω��RÀ�[y��N�xT�=��[G�jL�iW5�CVϓ�㒯-�e�r������˹��ma��ӦBW75�������9�dl�o���!�>қ$����Ǉ�;S��<�"g�m��?뼔���H��Q������7����6����'���sk|�n�o����6E?�(?�:<��TK)	'n"q���(����;�↖��`����v&怹�ݸ����@��f�U�͛G��z�F���~F{��O�RUo4^Z[^�e��!���|:/q��1�v�}ė�
��,`�H�_#��h�I�aU�����P<&�����I:M�o��_x�����By� x�Bd�&R.�?$K��9h��v�����Q<M�kg�\r�.�g_�m*��V�_���+b��p�b�bP?��{��N���Nն��&?��շd���X(,J����i�!,���X�[�8.]6�?#5��.?��@V� b���+0���&&&�ݯ�}肍��Ӆ�/L'/�,����j�{k���-�h������|
�?�����s����������98�Y��q��E{g�F��2{\�wD��ޖ�a�L}w<�����(!�ޛBR���;�W���3R!�؇�ñ�&��X!�����w�}�?�(��u^�9����`�3*2�@��S��6}��U�1SR�#?^\W��8ꖨ���~��yk8�����K�~nk����J$�*+�ӧH$�",q��v`af��ϟ?��E����6l�*B~Z�_Ý(�dez%p����*�ȇ	�k�C����1E�Ά7Ȥ�@���y�����_�����GN�7y�<��IQ��z���_���w�/�OZԎ�$U��(�%%#���K~��E��Dh�������ʦp*�b�c�t�W%J\F�y6��pO����Z�ڔ��J ����_�����)�� ��]vwt��ƥ6蠒_+Rp'���Gt��)���/c6H�N�a��`6��W

���3��[=߿��x������_���d���]��a�|1�G�ٓwg�q���C���"�z@�xMeE2�&x��K�(�`z�x��P��kt�5�l&~==�N���ź�����gƾZ�y�J~ڢ�g���h�
c�9S��W�6�8�7&A��g����<�?R��'cUWf�w�S����U�YxyѢ<6F�?� �G/�}�����R9�}��Ѳ����(@��]�Й"��TI̍��7�P��0}V�T�~8��C�����a����d~�]���YY���y��y���`}�����M�|��gcQJV-��='�yP�����j��;Z��>�a����	R�[�;4Y���%/M~�����dKxf�����wcD��`���E)��^��-�C.��S�ȷ����<E@):-�����V
G\U-�;�'�=��Z��D!,����QN	iizI�����S,��?,�mZs^�(���aS)*���~��i���?��3.�E\碟�u����
����0MV��+�؅�SU�f���?��6��V�{�RO�4��A���]7��L����������8;kiV�p�,;A�-�F�rp���!6��oibS��1�23�����ʓ�bF9^����Vn���ƍ9/Jf;XI�@QQq�/ �Po3>*�0��`�=n�777�ߣ٭H{�{JڔW�r�aװ1J�J]�6��1GG�I�Fru�J���1�S��c!��� =I�Wr*�x����SNhr�.���7l�^<jpY�9ށ�ևþ�I{?�^��Z�=���^o�0V�?��1���ݭ89��o�x��_;��rQ��ݵ�V3A<��x֌*aƆE=��7X���{���0OqG������g���+�?U��U����Z�z\^.s�݋T�x�\`
�[�#��J/��C�d�>���޻܀,�������C��-�����.5I��,����5����5���W���r��.ЋC�w�>��Sq�ϡ�-�;Z����z��>'<	ʖ����ߔh��&���̿B_C��.�.�v�žt=L����(0UU�U|ޫ��c�b���ﶗ��P~�ɲ).��mCG憄�4f���QNVۣs���Ɗ�nn��3�P��Y;�Y?!����9��J�&�0e[��}�C%�Fô�+� ��,.�OD&���@�nh����x�~(���m��4��'�(����s�h�%���z��3ظ�_�a��/�P����2gIn7���L�8�L�;R�`W1D8��Ow^�B�^ܥ{�������m��9�r7���]F�^�k[�������kRѩ'>���}t?=ݵ����������#rӖ��҄����˴U�#Q�Yg��ir��
B��5nLT�ޝ:�3��{C^�BAA���H�~�75��^���f'�Q_O���82�Tcp�ѣG���nS�R��5��c+�GY�����_���
�4��u�iK�i�5>�./���',��η��g<�y��x��#[�F03Li�Ԛ�q�i��SCv�#�IP�vx©���H�X>K�V���������~��H�fw�6��B�"nߩR-�]4"�u�s�&W>�!�z濶���%x��N��p�O㧑b$���$�Nuv�I����˅֗�/}zF�?�֍���#ٜ��q�k��u��]8�2�612�9=y%�R�EM�U�KM����#9 X�U��n����������D���FI�ذ����O���͍zO@A0��!E���JA\�W�5 8(X}�����v�V�Z�`�����l��Y��}cܭ�K����S5��HOƛ7��^3&l�Չ#�z<C��v"X	<�F���ng�{M�מr �����,��{��r����e�SL����C���8��)K�Ɋ[��N�h���q�r�U��������NʇG#U���O6����%�=����g ���g��2f���b:]���:e�,��˹�m�
k/�"b�D+�$�QL�������Ш2�_A4}g#d�0�=��uo�ex�����(9�A �c��c\Kۭ�����zᗝ��ve�%vޮM��ݬ���Iy�w#�����1aA��:!�3�Mu����#^mv�WV�jR�=�ْby�y�����JzŰ`����i�:l�'��
{ӓ��u�M�R(����׻�ύ�2b��g���,�3�`�m����p�7;�!�.5G�ns>m�H��1s�߳�J��&~C����{���3}�1Guаz)!T!
τ�gr������!��1���܀��@1�B����&)	����ܲ��~���=jN�YFo���c�V]��-�y�f*�.Ѹc�F�q�Q�S�G�I�����elj�=�}q�!IS�ݤ2@Y��M~	_��&]kn�mg1�O���$����d~��2�ޜ���J�Zi�js_-~4TZ�U�-?1]�{���{L���ü�a#��f\����;��o�*���CQ�F�8��:a��E Y�gAK���J���4�����Pw�z�NM�/��q�%\gD�^�I���=����\�_�`�n,�&�*>�HpΓc�ݰ!?2�{�����~�ߡǄ����	�#�v��/桉qwr�}S�>��J�G�cb��V���qT�P���|�`��"�%C�2{�d~c���'O�p>���\嫴�UE�����QI(�M�?�n�ɢ'���WV0O���S�c9	7�%���=��/n��̒��b�;��qrw/��Ö�3x�N�ñ8@�F�?H����T��F[�n�FW_w�v�]:${���Ku���'��8�dc�+��5�9h�w���e5BeUF>[�zS�������Um�0��/��n)6D��>��k�M��݅����r@���ʕ ��\ȠNj,q�Hś&���NU���W��RP�hǶ�{��6ez}�?��gC1���X��	���:~���"reI�K��(⒒��X�řъCZ����&�\Y8:^���9�8O�K���Ki�##�^�7��1��۰�Za�p��`9f�%dx�_�9��%��BP�@-��fZ�7��::ư���[H��>��gz�70z�Uk�:k;ɨ��۝�>�˿�u���1�fD3[�v8�ǋ�}����6�=M�|T
(���/���(M���E?p�{C��azQ����I��iM7+�i�c��/S�������~�:"��=ӋXl>RA��K+O�b-]�� �j�l�=Zl����b��n(`�	�1��t��ߧ蔘�����ﺯ�<I����-���U:�I�]KX+��ǿ�6��PA'���r�Ҡ1�a�����Y�O|v};-\~8�!c�1�,�U<�5�
۷	H3V�D��+����!!�&3`���ww��7ǭ)�%�zeN}���{���9�(��� �	��O.]-�9䖔�z���gg����/�QH��a]ӑH��a{�:�Oָjz�/ZS��5���D/ϣ��ͣ��"�p��PI�G�5��[����8�*x=�%f�:�Ъ�_sT n�!�Js��e�O��Ki�IJ&V�<��w4��m����^���7��N��"�d�m�����V___�2�塈V�$D"zK�xN��ꎳRk-[z��y�ԟ�ȁ1�=4�K|$�����.웳������W<�Ս�	���i�^��ؚNδ�aEV�ơ��6��u�#�\���T�d�S����BBB�#�x�S7����Z�Ѽ�f͞ �$7B�.���Y0k�a�������bm��rB����@�.4��h�=�/�?��k,�V;H@���U�����
�7�N���ro%��%oX��Ic"7�_��%�}s_
wLY_n'�ޘ���w�*����"��|��*lw6�����K2�s��$V�^g���{z�#��UtvN��a�����JN�I���'�<��rf���.Q{{��
��&<�W9��9kl�]K��@�|�MM����h,��Z����*�:!-��T:�]�^�����S:[u����%Pe��b_}-,Z*yV]!lnX�|�aC¸C��N3���u��89>�c�G��D�4A�Ͻ���YV�GSk�D�2Wq�3�֥���W�/�QGH8Ͻ)ؙ̧ۢ�A9�#��j��+�s��::�p33G�i��G4�S�,��|��qMбw�V��=ƍ������}�FshfGo�x�8ϣh����ll���
�k1+�8$���Q�w��B���!��� �D�H��y�}i�����������g�bn��I��dHg�G_���XEE��s]%8��C����*�:�ЦJ����K76�o�ݗ��qt|v0��E;rK��As�������X�õ�4�tpQ�\��H�2 _�8���ks�gr0���u��˛:���O�}� �Ǉ�h;�_��*&�|/r�?x��J��f�[�H�-�����]��J�s�9-ͪ��x�~aq�+�U�j*�ң�,H��Y�o�H��|��d�R /K��C��53��x�P�y�h�Ac\i��� 2GԹGp����G�ʺ��-�O8 ��h5�FFF"k%)��:& ��=�m�4�z��ٵ/���K�����w	8??*y�5g�d�6�@!�?ܒ`��a�¢������{k�r)B#|m���T��G>`���������X3��'~�͂�o½���I���lg��2h%��g�9J.zm%'�ĉ�.��A8G��ڿ,~��Ȋ�iMի�{̕s�^^��(�e]b���l؊�-l�M���q�ϟ?��<�Uxg�Bpǋe >�gr��O���cn�ݬ�Y���_����+~��<6ovg���}���y�`g�j�D�j2�Q�x�NN]�y��uZ,NAu���x��\ʎ7y��$(���L4.n���邺+̵l\��)���&��.b�D��p��W/,�I�
B�}b�e�˯��87�!7r>?7�K7i��dC>���鎙aE��_����q�!�]�a�֌��J��̜�_R
�k���]Jqn^e�q�ew�k�;��9��]�5�3p��a�%��ݐ�:^�s��꧖0���e�g�4:�afJ��.��^�0\k^�H�l�h3�H7�����y6h�y��6�m�6�����i��r�VGK褉bY��7�ꧣ�|��u.Bp?��	�~�m���<F���;L*!�$h�Wa�.BLXz<PS�)���|-o�R��OM�U����l�[	�<`c�J�}�~%=:�I���			�#�:#!�>ZP���Uڨ^���Y��=�#:d�9�~|��5�d��M�et�N/�|���spp���?T���bJ̼9�.Ƈ@�'������T%C����Iߏ��xg��7����Q)7X>_^����}��mKqv�߫]�e�+���-�m�ܪ�u��	|쩒�ߠ;=2�#�ڀUڇaT���at-S�IQ/&k]k���t���5�~߱)�OS?��������v���4c/B{�͝<'��ͷ��͙�q����Y��,�@��7��+��iZ�A�$m�����$��}.��(����4���ƎWYEE�o�@�A(��#%b�hl����\�����h?z�P����ߝab���B�br����G�h:yrN���"��r>��
L��s)�%3�]2�l�#q��[��7��u�C@
-a+2{�7�oF��F�T7[�(�J�*���^�D��&��w�[���98����F:7��'e�p�ʱ�Ҫ/�N|��&ʄ��$�Je�9�a%����|W~��%C4��j���Ŏ��,��}p�
��I�7�n���˜�G@�y��l� ��<��ߚ;����
昲M�^ڡϯWX�ήP�����e1m!�Bl¶?>����_ΰw����[M��5��#�qy�븷r\bY�t(�E6��}��Kh��tb�Cܼ�l�T�Q�S�l=E]ϽK�#Cv@�غ�վ�-ed�-wPy�)�\3{�l�C����	��������~ۚ��AGl����,�B�_oh�i�Mr�&+:���=9s++q��p_ޕ�>v��~rZv�&��Wܲ��'&&�k:z�5�[�f��v�������k\�9pYݑ)3�b.	Z2z�H�ol?
�8��M�9&�d�R-/E"�/�,�;1eB}���b����7����$�2֧ty�����^dY�Yo�_:�W5��XA�:*�|����T�M�V���i�%�1��H��&�AP_������ijxA��wG\�?0lns%>�N�H�G���^��X��چѓ|�T�H>�x�}�(��4߷�tX���F:U��=���X;���J"���?���qЉw���p�[<��o~!�n���+C~��t��ҟ�� =o���U騕�ö6�v=cc�5� U���ls"l��h��"1LK�)$�`��g���lGw��v0W��g�xP�4l�B�l�Z6��1�5���`��u���l�����|�yT�p�|&hZ�K����}���,�7�����m��$��A�<*o�8��P�N���L���y�_N�W�.�	pq�w�[ɾ��ҽ��u.��������ۯ�ڑ�V�����fsK7����و�s���+�[���5��|w+�Ȯ��0j5@�Mf��)����9�Q�<&M�D?>�-�'���{@Rb�	\s�ɺ0�ģC�c���	�R�A�o!.*د||�a��k&�F�������]�� %L�E ��˅��;�{q:�/~{�������Q\G �>�|��v�=9y�[�2c4mH!g^"�Z��y��q{?�1����R���}���o饒�0S ����?�97�g|j��0 �)6�PY���A0x�J��1�P��{=3s�^��Q�s�[b|�����7ox&ȼE.
Ժ�tB)"���m,rѯ])t�!	Pk;���o*��8���CCl<��"�r���,�tb�%�����ښ�QYU6�+�\��f��\J�pAh B�m�Ep�+3Ff���ww8���U6�@Q�x�&EF�)�+E���ս����b�o#Y��:�E �F!Gz���[��3��{����'U����;�Ahww���>o:F � r�5�A�JFK��X"h�6����Kl2-� �˛R�{w��T���ܦ4��pO�1k�SZ�y@[��
�6C���@�|�څ��ì
�����߫9�/P���/�GF�C���EFs1ՙ�����e�nvuuM�����9�#mc�����4�|	0�$��W��~�p�t+�;���.�cq �uʒ��r���6�^h**�hBSL�'g��ɦ�_*������4oTx6Z�Լ�~t�Ձ��1b���d�W�s'�ܪW�)r�렚̱4|(��m I0���zҠp
�oB����d�a0q�����}1�ۋ�����=	�,�S�Ճ���G�c��"h����M'���?k]{��E�T�۹>�Q�Or~�薔�e������� 7��"7��bȂ'���f@��k�e��p���DT�c��y����鮾���Uz��=\ ۄgqT�W"g��".֏�B2!L�@/e�)(R�n2�B��y�j���������,禧U>f�mx�ż�G����?7]e@�)�ߏ�"��r�'ռ�p�b���H:u09�'�Q�/�ң�m斘����+Ę�:'�~����k\���"G8)x7δ��k��r2R�*ҡ��2�?K[��byӯ0T2����pαC��<�&���H]EX�� ��Q j��N�ڨ���T���Ϸ7�ﵵ�Z+uP�`"��-�����M��t��U8<��c���ښ�w��1	�#2��u������?�F���!$@k�Oy�#��v�c�h�ƍ�����fR��Aǎ�}	���SvG����V?�X>L�,�����<Ah?ޖj6`�7�8[9��ǯ�%`|�vƀ��{�`$^5�����H��p*"�j����M��9����b�Ҵ������q۴%_9���P���*�"� �;^ai`l��xx:<��KK�LD<�h��%ݽ�˖DA9�en�G�@^R�F�T�ik�>���;�O�eX8ER0�fM��JR�k@9qD���1{Æ���2�5���?��yu��p���zW]X�x 3l#Z����#�[N�����`S	�;=
��H�#�dqVI�e��09G�,�/�r���k��Ɲ��ό�9�Zێ񘔣�u<���g.�J<4ֵ4kJM��a����6��V�trN�HJ�?}�pp�|?���E_�T�H�'��F� =^_���LMM��z�����K�6W0�����iK��/�
�)dF?_q@�|�*27k���E{��5*z���c!5*�e�͜hR�Q��,[{��ϸ���I�#:�<�)�0�I�����d���?C;(!}�H�SzZ�t)��w�����n&�=>���n�G��b�,����Mh�`h�O���x�"�[Y&t��[�����U���WJj�
���؀	a�(e�Y"H�`��)͉����iM�W�G�Q��ʓ�_#� Q�{DnsQ s��ډ�''%e���Y�qRL{��U?��L��E18YY�d�.����Q���Ãs0gՈ{�S�ޙ~<��~��O&V��w�Oz%???���P����h�Jr��O��� Gb`�"FJ"��8��0�9���U$Z'xh������W���<��Khk[��G;�J��I�Y��׀s]�s��~�֝�{�щ׏+�a�LJ�Vz'���u-�*{�6��a R�lڅ��ׁЏ��m��sp�����IM'�o)z�(!�����rS_�/�/�Zk@uoJ�uo��l���F��	\���lw^X��(Y���	���i�m����Yt�@��ˏ�1E�MU7����ͧ���i�=ĂIS��n[���iσ�F��Zzd՛&m��Uo@��n7���6��q���h-����������$%��e������(���o�#{�a�LT����%$��3ٗ���uE�q+����y�����[6� �5�S6-?�#��N�N�FFF��rH�:�tb}�qꖽ��2��ξN���$̮��y��F2N^�\L�2҄֫����S�Eykˀ�q�{�7vW��u��6���G7�yyuk��M�҉w��痋�>i�;��"0���pң@��4�ouu�����oS��m�ngg�},L���k0ZI19�/]7�E>�}h��h@��ÀHn��x���8���;�Z��[�7��拾�A�p
G��x9��7@�m)�O��aV�ƭԍ���\Gɦ�22�f�M�AL_ƢP�y	P�&���@�I]Z��@��1�O��mti��]�V_7����� �7��b�q�C�M1�[�5��.�(&=p�0)aȕx_H\��(u[ ����0�MO����49�I/�[Z�줻���Wۉޮ�?����o���3�6�^�|F@��%Ի�������Ζ����	�sg�1�pr~�F� ����箮�Q�>��h~�:�z�^��
�m�DX)7#�,�/��;^e?Z���p�C��,��g�G��'�ɇ��o�fӮ����[U���Y7�@:"�J%��[��y�4�JV�ݣ���a�I�M�������(z��Ǐonv��\���ꍰ�m�4��u�ro��~n��s>��lTxlL���iQ��5����R;�V��녺��Uܬwl��8"LtҖnz��~�3��P�2�nL|מ��F�X92��|�`c�5�����y�/�0��wKG�fB;d�;`dݠ�����0l[�D�9�Q�NЭX���b�oT��^RR�B�ɠ?W���{��?��;�F%��^|��x����J��a��-�Q
����ȋ��-�)��oc^~���zo�Kt����%r?[�J��A��:���k�!�[�G��]N���,C�ӵ��&�O��.M�N�L�Ǚ���y�!�������z�*	���~n+�]��_J�~�wX�߰��\�0�L��kp��Β��q�b��MX�c[�?�l��环�髴44L�C�-�@-������
@B����W�����ă��{9���}@�T�L�_��fh��芿hV�M}Eٱ%����D������O?s^$�9l����J?�4�N����o��KBL{��k���*?#��\���~���R|L�^����{�?g����ׯ_1?zz+;$��#Yq/�^���߿���j�T�+�ܷ0�o��_s��^�$"4�@����|N3���y�^������q�r�9~F19�>���N�ؾ@ګ-S7�]=�Zd���R<��= ��$�JI�����R����b��"���L2N8�~�lJ9�.V��a񉮶8TO�SG�%����8/1B�t���1����jU�7�bV/��q�r��پ�kZ����аR����u���80b�&?~��~Ex����Cd�r4�Q8�zZ���h��N�k�%n�R=��q<�/S��$�~af��`x%7�����&�0�|�2�&z�@��=�h,f���B�N>�����F��f1xؓ���c��MX5L��~��a�쵖�r��>�uP�|�p��đ��?�F���&M���Ԁ�ո�'I�_���8
}�T�Y�}}Md^��>�\C����Ι��ݗ�(,��=ϫ�~�"*߉<xr����c}��5�������1�~��6�1M�����s;�!��o~!�wBv��8���4N�Ԇ%��=@�uP�[��Q5���N9%N����9��\X\�����1�Y�V�'���t���F�OBz�gP��k�AE��E�$�?�K6&d�+�._2�Ӎa�c'�8���։��R��?�}�h�i?�v�3��跳�=�w���3+��=�	�؋iKW&E�Z��8�3��)���4oW�h��:���zg�k�e� )Rw�t�;����AZ�L셇ICl�ư��n�e�d��2�P~�je+7M���w��Ҁ�?�XE���
��fV�Υ�?� u���8�4A��g{�S���!r��V��)����
���j�]��c��\����ALJ_(�q�B"�<���8I�S�D��	sQ���[�^]��=�2Ģ,����I8��C!�n%��i��xt�qQ�ǡ��dU�)G�hR�{6pGPC#���O��\�?H�"���eH$�~&�)�i>3����'*�˂�����ᆝ�vz�a��/��^@Yl�����_}�GX��D���#�л���>��k�O���r��-�A�h$2�[��8������Xeg�9�yۨɇL�?�S�ޒ0�Α-���:_�,�> �s�CbE�fb�CP���[�,���3�.�I��T&���:��Y�0���j�Fc#��QwA�pC�BK����%�����+g�&��L�P���O���G�۰�Oe֐���h�WUQ���J��ҹ����I���v8����RRRƨ;N"M�_]�d �1W����l����
)���$�)��bDF�dT�c��M�G�HnR�
M�)���K��YW���V����}	1��mQt��2o�.NwYz�6K�E�0�]��׌����\���āz�TH{ﮍM/�,��b���F����PN]=��)���
;�4
�f�B�Ȏ�g���"��&�k�􄓮��yޘ�3ov3S0C�.�Z��Xu:yte<
1�}^n-�ʸG�d��T�a�Rm����'�ƾ�>JY���A��:�]�Ã��ģ�<#�U��fߙd`��D��߁�:������j33�_i�S���b��R� ���v�nܦ	ӕ���Ȱ��׿AuJ���O���C��5�t�g� �S��a������A+����n����Z0���1���q�a��ͯ_�m�¯m_h!jZy���h��>�v�Z���{S ���H������{���������h+�A"]j�����5����A����D_�Q�&WX�#|�y���e�)�?=9V`xxs�V�{%�YTL�9A�J�j�T���Щt���&�gU`0�6"ufK��y�-z�a�����W3����,,TŇ������h�ʐ4�9��E�)��,�T�$�A����(̈́Uf����&Ok0�܄ʼD������0\�ၡppF%�mn�����%ɉ���X�B־;N}���Ӊ�S<]������d��ZV2<L��NmI�@����^�'����Dܺ��u�	�)L8�'׭0$�@�^���}h�yTA�bA�5�c�U[
;qa��>3������:����Jz����ſ�f�%</e��ޭ�[�-N?9�t���7��FWN�v7L�%|������p��kɨ~�gϩkx!"��H���$V�ۅ��8��ʊ����4ܔ (��)�:��!n*M�	<*L}����l�,�Q&mb߽{�%!@��;�����,1���iv�l⿰HFݢ������
)����T�A�7Y7�ipΰ�.����!C�D1�Гk=v$k#�@z:@����s��E���PSni��*�I�d�"�_b����NH k�~p�����0J��:`0N�C�T
�����o�T<���/õ����É*�^_����aP�I$9��X�_ːUL�7���2 Rjjj���ޤ�$pe*�h��P#9����l�xk�>�FP��c�@�X�������)E�֎P� &�����<#+�ɕ�,�#�K�P'�c��a�_��������0�Bѽ~}}}ɪg�Z��V1o�7[[�b�%0�I�?�xhn��&������Im�`5@��P)spkO�	���?W�n.t�����hkLҷ��Jh޼�O���l�!��5/�6`��"d�\�Ŋ�"Ѯ@e��I�*��0W[�4!9���7d8��g]�Z� �2j�K�܂B"l%2T��A �o�y�
��W���j�P�V��MĎ<��"�p!��{��wT��p�C��Li=z�ͯ�ŕX4cQᦎ��L}��	pW4��*aCP�|��\�R!�Y?�����,Es��Ǟ�BO�Q7Pa��R�^�Oc+++�ѯ�b���g|��FZ�c3@�Mi��� ����z����&)���b�	��K��T������R�j�"~"���罃��������o�ңa.�XڻK�e.5�Eύ�B4H�����W�Y�1m'G��Ɉ�(+����]	�������A�鋸�Wd��}�l�N�|h�t�L���������;n؏�C�����J��Q
�*jj����v�!G��n�@L�����D����o�;���l�w�����������$矇8*vO_��g�M�7ȕ�s{h���B�*�Q,m`��s:��	$�͑�u���?��I��K�	&�����������N�P�@��P�Hl����ױ����6��5�k0P�/w���h��F��L"}���KB� "Yi��j�<��eAn��d?�A���d���	Pnؠ#֬��od=�1�B�����4��հ�Ka��a���	��ޛ&}���>�y�B�3i3H�Zh	n�M��o��%�ݿ{�h��RC[{���(u���cS�_���[�6�fՌ���;�6�Ҳ���,@��!�LiP�F��=�g �eR��6U]V�"*	�'uDU7�"7����"����Q;��q4��eF�����$�%H����Vҙ�"�l�Cf������Q ^+y�iw�>&;[ZZ���8�#YY��4��h.7����$�K�
��o���:zv�c�������v��%@�R��D*�Hc')��jkm��\V��d�iDu��p�jz�6 UA�S�L�	�d�������@#U��U Dz`�jA�34��J��KO߃8}�Œ��u��,:=1C6�@J�����S��	�y����ۇ_gf���zsN��y�['������ȉA���y��V�˴JPmm�KA>�,F��}���u�7�2ϣ�7��e��g ˌ�UIr����ך4�6��ԁ�Ӳ�M=*KoÇ0�	��`�8o����93���f�Px��P@�fᰊ����az�t�p����NpmW3�y�^%O,��I��cvcU��5�����d�J��]b^�[� z�Q1ۻS�;LZԘ��=�~���F�6^`�U�o�h���Ei��p�V�u�����x�!	�|�!��f��3O*��?��WT$�-�/"%������T#���)���X:T����c�+�ʣ᫪�Y�ձU� ���
)*	
W!�ydcgvVS�dEh�����c#	n-�M��9���.U�O�^ ^��e;�N�ڂ�ː6�� ү���V���!vs�r�aTGx�+c�=���ʬC���ݻw)�~ P7S�
ȗg��'w��
�|�#Ľ����m�� k�WىP� `Fԁ^�zk3���BJ�?�"�L�4�׎�Z��F�񭐿YSB;7߽=��@ZB��*�ъӲv7��ұa���� k��GW��5p���C�L����us��|`��k��j6p��Y�Q�����eƦud�ǔ�a � �J���{^�"����rk��K��<�:����r7���E���2;�X'���B���gV��w��7F݄�2@ �e�c'N�5Yg���f<�(��]�?���{؊�0 s"�f�K&�．DҞ��q/��$�_)���!A	Җ�Ux���]��3�-,,��C��˻RO��&9TaE�"̽eB=~��>����wi�?�&8������6����D�l3J�87Pz�4r���R����J�\l��?�&�| <*s�5���
|�G���p$7|!#�!|��˗k(�B�tگ���
ܽ�V��5���юX#�o���t&�Ҭx�}�6��"�P�D��>u�o`�%�P�xڡ"3��i��t�ߗ�ߛTd`�1G�2���
��/N�1�wi�=@��2��[��vgy\oD�j7+�-r���O���{c��̰�(w^�nB���"����z���wҖ:��|��
EYLǶwR�m{�/sd���=��S��ӧ`��0(�u=K/�k}��9�i��Ä���,�k�Q��.3�X�<�F�b��5��Bh��3h* /aҪ;��{�X����*�� �q�N�� i
0}Ǭ�{P�p�׊���k�^s$w��5��BC;ZZ�,��^��ajv�T����@��T��mwm��6��
@��U�(DK`OO����ӟ�0p�	��M�\�>l���+�s[�/��8���)��x����������
��b��R�k
d�K�%��C@X�����wwUH@���W*M5�s5�vs����kD5i��M�aQ�᭙ ��3�d2<���n|�B��\!�肿�[��z��ˮ����-Zy�����K�wp��������=���������)� U0�/�/ y�|�`:;n�nX���qU ��<hO~��9W��o��M��%���o���X=�@��������w��EU㹵�����l�(�]�G���sp��h�aK��*m�yܗ�H����"Y��-M��y%�\A��J�
{ޙ�Gw~�TT\����㡤�Lٯy��:rϵ���nacå!�����*���/�[!R=(ӕ@γ�	�c�Td�0\�uo��&*)�}@vh�����8��� ���J%4i��Ѣ#&Ϡ���ⱶ���Ťk,��b�\T��\Uݯ"��RzguoIy����Ѫz�Nv�9�(��V��.��v��-���.)(�?�%�W&1�9l���ێ�tYUQU�����n��4Z,.�ĕ}�<񎞟�~�Aqb/	���@ݵ�����'��!��K7d 2S�x������3a��g-d�%n몍�����=h"��u �6
��Io��ә�>���gk����@,ŧiFs�Q�]�38c� �Sh9f0�xtU!hߙj�.}�1�bP����l���j@����3�ۋ}Ċ�F5⎞�Q�$�n��=E����vKc���N���Y�S���@��೘.%U��*��
'�w`pVtb}�c}Bg_��,1ȁ^jw����r�1�5l��ָ�����	�PT*j�������/$PN���)e��3Z�=�O��Y���5<�^l�ȧ����?΅��0�gψr!�����7._�����Q7O���K��L��g*�}z�}vS�̓7J4��oM���QS��P7�HSS�!s�E8�{�1�K����_I��%�LE��!�j~���JJ����6H��j���dX������94��M�'�z�sN"��=7h��Ӟc�j��*��? 4]^^V�Z�����������������a�w:9$ ��H���ď8�S�`t�Ϡ�AݫR���&� ��z�$(c%������?����bׯ�u! �
�zƻ>Uѐ�o���� ;��4io��u���rm��L����۾� ������������0���L�%����xp�zV��Wl�����lm1�Z���'�:	���Gr�\��&�@9��Ĺ"�����
'���O�y
�pT_+mG^����~��3�d���J�z�$W"t�,������Q�ͼ�_S|8��sp���VIÁ�.�FpW�I1�΍7�{���z���F���P��m��TUU[�Zִs'xj�Ҽ،|�{��2P� s�����p&�1+�_+5?G:��߿W�;�>N��u��k�N��뭅�8�M��a�n�W��g;�]�_]�/+-%Gm ���i�1�sNZ� �?�9���$^"n�»*���̇@��F�F���H��Ƹ63]j�df%�y�'M`HW����B�7a|'�!�#�fl)��uw}��E�ϠʲהPSԈ�u��G�#��M_cjjj��_.�i>��Yd�*�����@�Q��I�� q+eB�j\�K�4M������o�g*��X�8y_�.|���0#v��g�KgF3��)�0��d����:lH���b��$!��i����z%�����+�ߝx�l�v�l����������ޒ�hx	����fy�<��+9~ ܜo9ݨ~o+Fda	gv��w3��.,�iװa%������{�p���xZ�)���HBY�,-��!�!K���(�=!�p!iȖ})�d;c��������}��z�{�����\g�8�j�|��~���k�?��0��3ݞ���:M�c1�ͪ�W�5U�`s�\'���Ó��� �L���N`V�Q��x�׿�93|'��,9��n�*@+���	���A��#��拞��FY�y����UȺ$%�Nf���>_{:�A���ؒ[�LBD�p�Z���ԝ�ԗސi�E�ۨm�)(�*qJb����IY'96�Ho��I���*�%U��U�WN�x�ϊ�~����L�^����[���,a?7������׆���}	%��9U��̬)�I+]��gzz:� ?C��+���vI[�A�_3��uzG��e����؟Ir!߃�/?����)K����e\sI�7�77]--��g��5s��pQ/?͆�՗���m�����>$�thg�˃���x��h��ǩ��������o�(/���m�m{���;Ix��֫]��!����?o����F.Kp骈5�[�cx/\�6#�^`���񫛟>���R���O�v,�
d	7+�=�Ƨ_�XL��P�Y��v�����	ξ�Q�=��͉B�q���מ��ݲa^	2j�ǉbT��f�tP����5S{���e�y�@���Q�]��}̸�{_]��y���n���'����|����'w<��c{u�yx�iYD_���***FS�0E�����ֻ�+ٌ��8I��ғ<��}�c><�7_"��%3d&=��t�"Ҏ�Z:lǒ���ʤ���%x�|�Bt�gwh=�h��v�i�Sj�n �E��]]U����I��f��>9�<OL�V���o=8� �]׺��>������Y������F�����J**�E�%YY�&''?�_�v��Bbu��=��¿�<���/_�������4�T�ͭBۛ���-Ky-w������u�M�eq���KmD=�>:��:�O�|f{Mi{ˎ8	L���wz|�|�1�h�$o
�N����k<ZW�8�����x�k���tͤ��"��x�O$%��)��/�\?T����<�ȝ@6H�̗�~���h��i�g�K��r
W�'� 
�Q�� uhl��@��w}mޣ�J:~�����~����$��%>j�䉎����y�P! [������K�OҮ[�tq't��z�������=d���}�0>����fj����A��B�z#a�ħ��3T�8�������M���%	$��yo��M�Ŭ��
��>�ΰ���{�(��i,��~bD �J�Vɢ/\�1�{7�S(E�f��q��H��M��W��Ǔ�EX�$��p5x�-�/�(�ο�hO�N"��|Q�/�.3в��Y-��ć��i�x6wS�j�.�7	���~¿���:�$�@�'DLd���q���x����V�����kegOz?�]�5����Pk�$O綳��b�[�N_�}�,��%(S�4�����I�������Uފ�92_�l3Ց_T����u����OO"�L#�b/j�512�z��0�iN'8�2�dO�tR�ߨu��N`���;^ �4+#E8��ą--9�ܽ۝E�hK�_kQ"E��#��Ρ������KR�V��d�g��� ���޿�cs}�ky��/v�b*bL�W�׎�����ʸ9:YwnS�*/z"�~5��u���^��Z�բ\`����-������<K�oPZߌ�jN�ˋ��R&����UPo9�ӽD���G�s-�$��_;�C�����E�p��2eh����`�We��x���L���h�5��pV��e�CI��d���'_�.*�Y�Ծ_������I롣�܋��/$��kdX,J�=�5��/boE�г�"�<�ku�Rb4�׬O���O�ꘋٔ�̵oB<���d�vp�3ag��}r�g�H�:::��U�� �y�+�b�3z�?BO�ٷ6 ���������ϯ�z�'Z�u�mc|�ܕ�N��xX�fq0��Ys|Ul���������rs�r���{(�)��\_h�ِ(�8�K��$��cy �&�-�cN\��ٳ�s���z�	גw�Ђ�*|a[�J͝�<]�.2�����|�un��c���v��U���^���z���w��+��$_�������l#��޹s�Ϳ�(�G]]c�2u�g�ڣ,<��BG�u���寖��*�/�a�a�puO�z���.f��Ƒ�m�'�ђ3�#&P�/���G�-[��B{���O`��!�/�=r	�
`)^��xf�/@+aX0`�.�z1º�Ƥ����f�lIX���GF`->���a�OB?9��� i
۽�~d�}s�`���<nɘc���g}&��@��(��b��O�����ώ|�౔n8���\����m�.,<�h�z�)C�=�:�<��E���D�|��مcm�Ш@92��A)�&�R?��ֺ�|"TJc��`V�⾄��6mÈ@&���Q�����-���ڔ(� D����-����G(�ǓJj\��Ɯ��٬Ah�"�?����.Nz]����W��'�����$��gP���>��+���gQ*%��t_�k�;�Z��\}f﹯�d�����2ɟś�e�����	+��+s�5���	�U�|� �p�ٟ8,YP]��i`sw7���u-��to^.LMI	���l����������P�'|i ��;�?h��o_���㗖��p./o���'̩<�'�6��굍]:.-,!�h}��6g̘���A����ui�Yqb��e1l��;����.�9�������n��?�^�����GW�Ǩ�3�;������R\�L�-�X�.���?��Z�~�#K����
+�w�5A�[���s�b�ѹ������e�TF���Cs�C-��'�F�[E����Ҳ��_}W���ằ:j��*��i�[�Ť�%���|����6=���sd2a�kJ2�u	��(¶rIE)%�=>�;��O��]i���]����׺Ҵs�����m��	O.Υ�z~/Ӡ��SYr�u.�?����9�suN{{UH���G�{y��M�̀3t�^]�/g-�o�9Ñ��h�[�9x�B+�¥>��J[�ku��u����˨q�l�
����oѭ龖$�|���M.NE�)A��\k�՜u]]��R�#��Nt�H���ȸ2?[IW��]3X$||�CD�e��lO��C�y�IE��@{�7a���'t��)�#���*T�#bԟ� 'q_�v
�R���o�p(�#��R"�u?G+��gt��'P�����o�n9��w.�bB��,����?ݵP(n��W����];\E����UOv�=�jL�ŝ5�W�����E�)�M;x/�_���Oy�D�7�W˰f`��y�:\�O:|pw� �s��L~�Z�y�"f$����<~����θ/Oɟ� �{��^wR&��&n�1�g��DQ��?އ8�%�����w��R4����_���0ʄ�N�q��<P?��C7*B�La��]&�7���Z��=��3+ncD�+�2/~��C�����p�7�+�V����}}^Fa�j*t�� ̬����&!�2X�B��G;��q/�U������\ƃ��ˉ�K����ɶ�3�2���a��ʈ��<DU�M��.xn���9I�����i��)
�vگ���k���v�d�{E�%3n��E����%��JJ<>�Z�c��սI8*�s��{� �~Ww2E�B�\^���i'Y�\��L�k��6ٞ�J��g�S�<�۽�z��f �BR�?n=X��dX򈡦%I.��:U=P��@���2д���9�%�C��D�ob$P�$W��q&x���a��rDM���{O��i��y4��r���6���P|s+]l � Ag�ROptvt�z�$w rE��pɥ�ta���%&��bg�?L<ѣ$츢ᕨ���0�R掁������~��ؚ��ռ�o��ٯ�̕���ޒS>�������dB]��h�������t7��Ç7;y��{�i�f+v��w.lxstik����öy����Hx�����Z������Ǐ��1 �y���V�;����8��~!B!��Z�i�X��7,�tO�ۮC������r��Z��2Ȩm?�����r�ps�Lވ�8Y�x{��hG]�D�@����|�'�
���9�955դ9^���c���KRRR3���gb'��[<w�D^_����ZO�o�;n{9I�}0D��D���������M�_lV���u�G�} ;N�&0z���}Λ�+�_hؕ������Epy�F���N��O��8-� I��K�$��ꪫ��w?=��?�����`�pn��kg���ov�k$?�V���?�סП�aE�]�r��ٚ�9-�� �XFg�3Ort��Fdd�l����aFY+��a��JO��{�,�˟<Y
� U��mDք���_��]f�Q;�ɰ�qaO���66(��z��F1G�0#P�Q�9b�79��!$*)+Slm��p�w_��^W�IF��OO��]�|�q_6x�6�L�)잷_�^��U���Pb�|wkZ�O�ٞTztwO#��+���_oy^��L��b��f`]��zo�V
���Fi����d��aP��TjwЉ�2�L�>Q���������C��MV���eB�v%N�"x�槮`�6��Q�51�!��Qg9���m��AQu�y��u�Ľ�ս`��m��P��q��:���0à�'N�˩|k���p�.Nڋ��C��[g��:�mٗ�q*���P�A멮3��F�^km>�2^�6ִ����;�]��bzۉ���wV���o��)V�1�)P|�A:�Yo)/�o�C��U��kP�S��{K�?��~O3gK�pZi[����&ҁֽ��h�%y�޽�������>�|kk��H��?�3�㛶��A�x�{��N�������?��Ν�*]p���:?y��7�:������ֳ�ޗ��?�D��/�[k���w��># ؑehy!�O?�җN1���y[�U��"��2�Y�X��r�|H��{��M�A�|r����d~i�B�]JQ̸�%����b��m��Z���.�X�e,^a^�Ҙy{���O�Y��/Dh��*JN/8=����+�Z�频�9o�����:E� �mF�/=�����~հ�bA�䞧��L����J���]f�q̕�֗�'4�By���n��m�~?�Wj�oM(cE�*����x���A����5��[i�O����1c����ʭ�Q��1�a�v��i��4���p�aS.��÷��ټ B�)��(��ǔ��nJv	ey'�6W�6WT�7{�	�FFLߙ����� ��ļ�:~�k��B������m+3�DOB����e$%�#�%R�w`^��8>/����2?TwWJ+�՟S���SVn.c��0� z6��݌���c� =N&^���Չ�(��!�3/�5�ׁ�>i������O�ś3��6xeԪ����'������ޘ. U����**��0�-y�,ll1^O"L�z����\.��n������ ���1p�̬,���(�?,�t!���\�LiZ�[iA<$ac1U���MS���:NKp}7��re���t᧼��0��ʊKJc�G%��� X�̒��Nk�+��,#�d���l^C7��(M��a"���̐fa��}x���C�1/�wuɕ��@���%�TR&�ccc�r(V)4~I��rs��ByS�24i�bG\r�s�4�9*EW��)�/v&��ǌ6'Դ���3 �H�N�)	28j^Dy��e?V�ɾf���VZ�0ڔ��_Y_h6+j\�pMY1&�	l���aaL���t&�}r���hPRRw���rg"� :� ���m���1#i�7йϕ�J\��K����B9�e蝉}�I!�w��n��r��˗g��4���,����W�ǔfӋ��aU�	^'��$��݄�y���K��%�*��(&�0�����/|��."���̥��7~��zT���V�i��v����L�b�?h&E�Tʏ60i�{�������$�w[KK�9Ȗ|�{�)�����:���x,�-�L�x�:pA}%q������6����1�1񥘖w)����O�u/�!�����"�pUrp�
x�ƨ���?���v[e+'�S�̏���D�c7C�:�?���w+�Z_d�tނ�	���*�}q�һ���>5�ʖWVƆ]K�Z4Iҥ|[t�xK���<�D����
n.镻N�ࣉ�W��i��V)�T	�H�du�aZ�7~Ah�9Xv}}T**�򻁕���d��@��7�4�̔�4W�c��a�׸𡻧'�<�&CMM�>h���BF��K?-]:�w6/BbV� ��qd�����"/$p���	70��:�Y�ٗB�j�:G�;��Q��0���@���7�ď�����vhH�˳�DA��|��i=�,��Y�7e-�$�'���o�^����9��쐀���;t�AN89;��O57�Y�L��x���H:��pY�mF!��ڎqQ�=�5�,�f)T��~����`蹤�1���̀��ŧ�������6�G��:�T�8%)��+���e��,�---UZ�232���f�7 �"m�ي����p.�Crs}�e�BR-5����� `F$dE�ɇ��J��ܠ@+W���J�P� ��h����<a�V��0��S1k��1GH���:� >�)��i6צm(��j���9~$ޤ���!���l���|��_�~���,��b�\l9��~�Gx7ת�N*/�����\J�d$u*��V��W �Z�]���sc-I��C����	�˜�u=(K��:��'�Rܼ�FO�b0��li0.7aR�5�\�T'�a��)�E�4������K�̞��M��l���#dE�,����Oh�DDD�\�	��1�����s�PK�yhJ��&�����ƕ��̦��� Ω������V�$2 N5�J1_��
�"�H	z?�5�zR�f����P��o�v��U.������|��$y*G���k����/]�g�M\����2�l����	G����,vc+�#E��S=��>;����_�����|X����0Na�� ��2��M�k/���_���;U�c�[ǫz���=�Z�P/�܉�ǵj�[����G?��]�����je_-~s�������	HU�L��15@���?�F��O �RȤA��f����K����̂fL�i�G]�@�Jڠ�U�Ӎ[{�@�g�K���qRk}�D���L��TR�~���2�y�??%�_�`k+����g �VC�)�	~�O=�$��L2��g�6�I��t܅��x��F���]ggg���O7�>�p~���+�Ƣ�%rxU�(B^s���8���X�cfgm-�e�ga�����Ds��q�xC,+`��A~^���Ƚ��bi�S���u@�ц�mU�Z�J��jx�ԯ9���
&|̖�0|R��0J� �e�����67i�y�Ns�r�I$�|�TH3�hⴒ����3��B|w%�|-}e,)dDd�C�X
I��v��#��Wi����к��������v{`�Y*84�8�����ec������㮏��8�_7ӹ{7�p}�)++�b҄�r~w�� ���[��R-���P]����r_��u�����j��\	�\	�
w����r����H�c�ۨ��2��JXⲃ|9~۩*����;��1_�Q�0]����pi}I���b�u_	Z�C�pnq�U#�x�C�UR��h*��@��X�&2�����B�y��?b}�6��/���/��v`
nq��>������p�\��3Q���=_�@B������@ ql08�8�i�14tl�1)���s��?��P@ZҪP��ϓԻ2��<��	?�U�$�S��u��KŮ�Q��&ǁ�4�k�ڽ���0 ����V�m��R���W㥰l�i����B8� ���d���9Z�x�m��J�ˇI'�����`���#����m�*
q_!�oe���e����7&��|,9_oN��:n �5�)/D��o6e���Q\�t;(��?�r�{�UZ���۟Q���{��zF��u�#�H��a��ؔSDf i&���$=��UW��L?Ǒ���2����+>xd�B�,PN��_.L,�iP����cR4Ji0&�@��	��/�.�e�1v-�;�V���ճ�j��o��C6כ7���	!0����
�W��#g3��E(m@C�{�������EYdS[��jL�f�D���Q:��
�0O�--m�S�/�c�����]�2�+5R/Q���4yl��J�d�)��bY��l^c3�Q�/�Bʃ ��~���=�z��w�J��N�� �rp����E���\uc�ڋ���y"
_�s��I���&d3hV�B���@_�;�a+++%�o�9�&���9�Z����q��d��ef8�Y��	�I�JW��H�58�se-���}�؝���l�J`�J`�;ɚ�Q��,�b�p ��sQ�y�����.�c-����� 2�g�&%�9/Ĕr:�Nv�a*d7��b*δ[��Vn�W�s1I�-�ׂ�qI������VGb���q��������	`;���%�0N`+�t�N��L�\W�Ҭ;innN�����RNjyX���t��
%�����VR�)? !���-� |�q��Ѻ��M�@�)�"y0)���A�IՓK���C�R�Xm>�'�)o?�����afc��|4�@D�/\���:`Y���Y�ٝV��؍���N��r��Ŕ$@]��+ ��I�_E��py�V�*/�f��s��؝F�y�R�B�ǥ���t.��)l�!@c�����B�/⿘�&�; �&� �cG_��u>3��o������O���Z� ��=�ih(A`�@����:�kU�������J$Ջ�]/�o78`�[4�K�������0)�2j�?}Az��X������3�$��LMO3o���L�]�m�
		ܠ�3����VR]\;�y�����ʀ�{x��%�t��J�2���{�{*�\�ҏ�V��Be����^��5�rv44?�n%˼�*kO*?��8H��j^(p]0-��
��>�u"�E&�Q�s+#.���&���=���i'�9i�@�]\]��@fwtu �b��Z���>�,����]��n�P1t&� �S �=X�\��H��?b�b�G��㳒�g���p�PӉ�)5���I�K�O�Ĥ�on�L3z�����M�~|����Ni��!���nyг.���u4n�߇n1���:��W��7�GHL�G����\v��a��!Prrrj�&�̯d�x�=�<Zש���#���I�D�ۜ�Gq/�j��d& =K��>]��ϒ��J:(-����/;��}�d�*��[�ϐ��l�¦0�䶦�TV�=����n��T��Ӣϟ�n%4 �lliy~�Dj��~3_���e�zX9��ұg�M�V��`�^��� M�h0�����ׯ��M
m-���D "�!
��-�s�J�8]--��6�¿Lo@�|_�z9�h�8���w���o�Mt�9d<�(������F(��	O��E2�6���=d�1L��#Z=��ׯ���	��'m��ǩ�}ț�͑�=��ߟ��'W���*�naD���~�����,ڄ�������ʂ���H:��egg��RHζ�8���)���HT��;m Ē y�/�'��Ԝm�^ȟh�  ���,�ײS����=w��q�x�F+�E�]��l�4��D?���3����@!e�����-���|zzy��'1	Y��P�����;�n��ipVSUN���l��8�>��ͳ���`��y��~�m�53�J6U���-�WŶ�ذ�V�4�� k�,5'H�\u���Fҽ>�� ��W�$���;­U�y�d
�c����p���c���Ebg<�F���v��;��G��P�@�M��P!A�HOu^w!ȿ���5Q��GKA� v�qFw��~�>�va=��4==N�|v�R�4����=��	���%�7�ίF9m�܀����L����6s�s���5Rvhs���0��s*F+FsD�e�.o��,4�����L��L����Wz����ꑑ����Vއ���Ģŏ�dT�e���{��$�Af��JE��$z��^Q�%�auxW����蠤+�;�a�z{�����m�����������ZY[W_%�����x�Z�磸ϐ��ڃ>��s��p'��|�?��߿�@E >^iD�MVN����uq9����/������6(����1�m[k��$!+��W�׋Q��L"N�fq����e��هg� ��r��]��0��]���S/)�a��7��t����h�G��A.1�@���FZZ��$pl���?�2�$�Oog�5���ww2NdT$�х��<�.�������4�i���y��t�
���v�]h�	\�y󏭅H���Y]�A�p%x0$x��#���!��6�.�xIϵ��?Ӝ� i�`
4����s�՘�qO��@�Ij�?���MQ��ޗ5:���K|�d�7�$kYHV�t�q�7 tP
*wz&��J���}]�}�X���M���T�%��ѹ����)�1������I5F�E�3�/c��}�xӦO��|z�ɝ�L�����&ϘƔ�N�0��O�@�1�&Hƭ�T��) �ׅH�1��ԅvʘ@3L@@M{�ݻ§!��ff���lE2�IZ������i��_�ڊ���+�!�t<�;Ԥs%KN8��r�
Z4�n>�*��ֆ,�%����ַ]ls�y@@2jJ�sH-�@Y��E�%�����)�; �s���"7�!�;�!g�����<
�=}"�Z�G�t�Y�y݂GIݟ��o�E0��C��;::� 'cJFϖķ������=��JcO�n� �A�L?�z��n;���}چ;MtqZ� [���[S�3n.�+s���Id�F%1�eђ:����M�d�<a�0��6�	t�4�}�˖}��4�i9����� �&:*���<I��Di$���I�H��Vvtw�ұS=$�T0���u�Jz[@6o�M}ٛzPa=�ĤC�a��=k��H$���d�s��ZyTϘ�Gd�V����r5���+�~ ]�}:�/[���O�l�bY�ģ���G�X�=�e���M��JL���!j�m�����^/A�#��Y�b����A1�w�����6�6��#��q���K�"�- -��3#۲�h�%�vvc��f�9"�ǒ%y�<f�(��@�fg�T�qs�4�lb���g����1㕙�W�ܱ1^ G�����DdT�P��L�&���F��}7��=@J�%�G���4\�96Ɲ�˜y���lk/h��O�ʕ ���o��N�o333?��r(����Jz�g��T����ʣ3ʭ�r������ڊ�٥���J#Cn��y%}"#
DK����Pp�����?I��ʭv	��m��[h�Z��EcC��?5m-�N JI¯�7�ݖ�u!�4,�s�E�xt�0�R
��@�|ݥ+�&:/�� �;�d�ۊ^��%�;�j-����]����Ro��[��T(�}y"�'��t"�}��{*++A��D7��*�����%rmQ�������^k�7C�J���2a�h�H�%*$Yl��:n��M�+ze�9xm2�Ɔ�T���݅������ѥ�����B�����N'㙃���7K�SI�r��c���a_6�M��n��K�>��^]�ƿW���s��xq_q����%q�5 0D��=�?��~�q�j4��m;���(�#;��m�|�.ݽ{Wc�:�o%�?��:"d� ?2os��U�-ζL$^�S�U�
������/�f�x30�K���ޮMj�S���J�"���!�ӊ�@�z1%Cpz��r��?��p�31݄8�@���J�DZ�c�G��Vve���p:<7���[S�cCu����=�ۚA�ȣ���S�&��~V� ����7E��5��O�r񇭕�3R��Kś�������$
;�GL#~+�a"�32;+ |P}WI.ӹ�7��?0����������f8�O����(x��p�m=MTLl��M����3���?k�;We����>�i�&J�^�fT%�^�z�Y��U)I�m�x�Ʃ�ӂJ�wk|��n�3���j�^@�We�yLYn��Pw@�˰bg�ڨ�� ��� ;y��1JѨ�v�[�C��;
�/�`p+E�r
2����Z��/
§��>�#8��d�Y���SCM嘆��?�������/k
��چ�X�u�l&�c�֩e2ET\<hpp0:���<��cAΞ|.j����l����1�ʶ�ķ���ȅ�oS���Lo�x��wB<���[��D>𿆔�g�F]�uw�^�􇎴���Ȱ���8\�Ӊ_�{2��1
�o�� �&�kdD����5�:�蹹�S��9������������6�z����tH����������@n�xeR��kY�M��w�a0�.R�cHy��}��򎀇;Kb����?V�5���=9X<���2����P�:V ��}�m(����w�ɽ�r�&���J�(�du������+���:,(�P@S󘦡>�_�	H�~;�$|��pZ�)$t+ʛȼ��s~�ُ	�:���q�JHC�0�b���� ����F���*ٲ�7��o�6
si����	�|(g � ꡧ�O�g?� )N>�{�)��'<�c# ��e�MI;0�thm!���Bh����X�'�1@��2\8�L�hH���V*�w��..��	>���,�=_��owo΅��{/�}�maA�����n:\�qG&��;[�pLP�e�>���]���o�" ��=�0�J��֪a�P�o�aBQ�i��qa-l`���i|��:7U�r��O��Ĭ��BF��YRO��5�v�
�NH�%M���ځq����v��qߎ��Y�#+6jJ�r���nT��T9�%�����[Ȃ+y(**�S��V���ϟM�m���T����9m`��%Xʅ�`T���� � n���:������3 5*M�g@6C�_
��HE���.wY�<2�=n|ٰfsc�BFh_~���D]��N
LP\½m?*�033�?�8ĥ�b9QJ�+�_R��V4>^j_LK�r"��>5m����2vvv6%��>9��z �Ҵ8��7��c+�v�\�W������I@���]V��)Ny�6s�{�RV?̐���Ve�#�4?��O�٣� >2`�Hl����rϔ�����S��۽�{O�F�Y��m7v��6b�))����XJ���i�����[^/�h㴌���?�M�ފ��r���}�+�l�!D���o�3�(�h��$�|���b�8��"��3�/z���a�P�Cr��I]a��S@��8-�+�A1u/M�V����a�NyHŨ((/ר�
�-�މ	4+(,,��
ݭO��v	XO��2:�J?�~�]��/��^- �vM�n��V���7kz� Sp \�P�#��c^���Vut�����Ɇ���<;�p����˹Y�K{�?�	G_J��m�L�X��j�f����<H����4SG�A'`iS���a��ɊD�X`�Q�ݿ��C�����jc��ذ�|�Ky��9�0�9�Ey ���P�(qPuu@��/ܡ�������n:�N�~�����zi3�g{6nď�Q���D�,�QO�=�	h��V-�1��g���bH|/o�0���QW�\���=��]���JP�і�贊��&�/� $�sr�2�	܇l�i)��`�Y@�	�jD�i3��}&���C�C=���s����)M����W���`�^�E#�P�=�i
�B��r���Hd;[�C 0AƏ�8,�/�h����֣z���h}š+�($s��bl����Dp˜i�=@KK����Sz���6z�3�S�0�Pκ�m�~�[I�]��FŽl��hu~eE�E寒��g�����!��l�ν�H�/�P/�v��[`ER��$*�kF'���W�<��A�u�Ng�&�7uw��Д�E_��i-��8�cRh0Aj���1�8ф[���#�j��N�M.�����Z����sT4�.+H?{u�BlO����U��-N���1=!�������
[ѷL��BGWW�wµ�{B��Y�}ֳ��#��s4 �sG1�� ����7��14��  k�&_d˦N���^jO*�i@����=�:���+ i2O-���By]�MS%�3�+�CC֏q���,�����?M���5��X,�I�{,"��L'�㽗z��aXf$���u@?������ُ=���H��Q�����O^�:������aU�"a���O;�E�d��d�����g�A�@�!`�t�/��>��B+j)C(t&:�u^w��OQ�~'O7�S���̬/�l;�y
�=�8���TH�}b��Rk�?�P{���]E=&eV�{v���N����p�H�\�f|���	��yK�㽋o?'#�ٟ��Vn.#�(D�)"�R>T�h'���Cי=��s_o��
�ޮ�?�S�f��g��yO �lll��F�x�zS���㷇����<�#��������G��Ӥ��V u1q�ۨ� 
'�?��1vр�qp 
C�F-0��*hO����T����u�+�s�S�f3���H���P�u:u���wh�����~M}(�I=&E���V����EYd�o*$_�Ny���j.M��8!ZHdP�(�
n ����[?��u����FS�y��� ��vEP@��MĈ[�_�+?�l�o�ֳG���1�R��Q1o��o�0N�񻴱��2�����=kԏ�ɁJ��m��������!@`��+��v��o�nr���0ۆ:� �|�k���oXh�2�+�a���hG�H�du�EX�Kn�0��e�V�����S�}=_o�w�`�����z^��}��]:<
0k�;]9��s�~���`ȧ�#�����0~L�.uwnɨ��g�a����zT%�3%���G8��r���������?����Y���j�5
�?�����k���r�����;��;{�cd��Տ�[��A��][�z�}5�P�����%j
*�q���_���(�A3r�D���l��p��'t��B���w¼m�\��������ͻ"�h�+p�_��N��o���-�'(dm^d��$q���N��R�a��g�^L��ټ��n�kj���0�F|t��hwK�[�������O�6�m6�m�"D�w���z��u�:�^O�����ީ=;�矟����w���>�+�>�@	��
����B��h'��M�u������M����hgzKQ���ݘ��.h[��HXWs�_�;���(���y�ȩ�c�߹�$���ѧ�W������iJ}y??��5{�f�k��x����5�Nm�Y^l:�6Hz��x��T�c�C���uW�~s����kѺ�u�Lյ�5��0���]㏬�T���X��ŝO�ݝ����W������V��[S˶����1���9�=}O�Rc�x�͍ᚐфg[�˗/��\z_J��y�����~>k�f/��8�a�<?ߛ�^ӷSћ��;p� �9m+5��]��jt'��Y�.������e�m�R��v�֫N#Q��!�����E��nR��f���������@0����C�����=מ�o���8X���૓�5�_��5�_��5�_��o�yʏ�칆����������������x�>�{sH���C[Wk(|ˆ�gj�ѿ���# ���*��g�)4{m�����m�fd%��z9
�T�����ݢ۬�?E{��w3�)4�z?��[����Ƿ�n�y��~��:Ro�QԖ_Vqc��r�"��ջ�}�/X���sU��O�S[�}3H���L�w��uUY�!T�4��������
�O%���2*�7�=�� PK   �e�X����H   C   /   images/8e6e9996-4250-48fd-a42c-980e5b13088a.pngC �߉PNG

   IHDR   d   4   |l��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��|yx����=[2�=dOHB6H���Ȧ�
����R��jk{�t���zi۷������R�*b�V@TY!@����=��d��=�L&$di����I~�[���g��9Ϡ�Y�����b�x�Ǉ���'NwC�R�j.�s��u�B��Z�?q�'-jJj��c��c¡�v9�v�w,��G�O{5:L�	}xߋ�mgI34�o��RB��h-��%C����v��:as�q5��Q89O�2{{Z|؟����,{r��
�:6B�U������B̞1}�������N���*�Z��Mya�������\.}2��Á��V��P+ZL�o5M`�����3�)++3(o۾� ={�ɖ�j,tOrL�_�:��E�]�����������S�qy��Mʰ:7�-Σ	��my.�cA�	Ĭ��Q�Oar�e^�3<C��Y�e��w���k�5|���Pw-��X�'V翐�����mGOgZ�.��e����@�� B�@t�Q�֪eR6��f�賸au)}~\���e��^\���RM�����FNz2�:��i'���G���E+�AH �F�9D��59�X��5;e��DJ�V*����8~z�ɷ&'�{%8P�����V6w@�V*���j4t<5!6�ʖ^�4t�	Wx\HU� c�MN����H��BhH04�h��h�Z��׏��v�jơ�N�t�`�0|=0,�H�����c0(*�I�t@���p{!���1==�s�0-k<�b���@Q@���fC���ӭ�8^݂/��Q�a�٥5�"96�/k���7O�}s[��*��,�AV豿��������7�"�X[�������i!��T�wAI㓑7m*V,�A�ށ�GK�i%���p��Ac������D�.h�k�W�I����~�(��f�c�iț<������zss�`�utuu�HI����k���U���� �m���Q�D������*�
n��Wb�j�3�
��	hii��`�
!�������T���a���������CxsW��c��'�e�A�ų"`�*Fŧ�jZpOON�����W"V>/y�%!xx��#8�h)���D{{;��܌��^!:�����0aRRRI�187%%a��|��{��8��.�O��9��zΚ��-�I6���+������������ݻ�u�V�<yR�Ɏ�d�J�PZHFF�.]�U�V!++	I����k�?�8�����e�U�5Rg�w7Y�ƣ��	�"'#���?�>���
M&�yY�F�҅�����~I��r~pЌ#G�࣏>�W_}%��K��S	�������E��zsss1.:wݴy�����wa{�����I�ya0R¼x��B,_�� X�"�oߎW_}� 5�e��F=:G��Y,�8q���X�~=��<��Cb=�����"�����r�Pغ�f^��һ1))ڀK�C����}&|Yg@u�Opc#X��S7��{�,CHX�X;�?�	��n���3�*��+��y}�x���
Q�w�yG@�я~���Lg*��X$��ފGڅ���9���T<YƳ�Q��Y"q�������q�F�8�d�PrK� MVE���dF?i�iP����_��_�w���ϟ�I�&�?P��ڇ�]k�83g-2���Rf���$���g)�C.L�g�ñ�%y�B4�9ߣvS�䖟X���X)q�l6�7���/��Ʉ Zg�&�ؙ��
^/���t�J�`��[��o�>��7��ʕ+����_~�k�-��q6&�&�f���ibFSS~������iub��� L�LG�����F&Ǉ�h���@{[�O���|�V�Eyy9x����X�b2H{��ף�孨��H�c0��`4ۄy�"#)
��:8u�A+ٍ͋9�0c�x�t�CK|>6"�m��n��¼t4wP\݊�-2�G�����߂x�n�Y8��r��100�g�y���D��`�൦f�#�,��(��C`��Bz��q���vY�^�Ǐ�cqs=� b���Խˡ7��%6ӛ
�(f\+��������i30uz��G1�?%��9-@�]\,�f��T)�ع��� �F#�q����Ǵi����v<��ð�Ւf���z�"��ff�AO���!� ���us�VbޔT��eAv2��}�
'cJZJj�x`�l�,vܺx�\s��E��?�Q���o]���q��>��h7��C��&�!o�L�Q�~v��1�x ���D\�R���܂S�J`"p���{N�����GJ�<~�BԾ����HLF��G*��U� <"2;v/~0xL��M$���?�ȄU�O9����Y�/Qdm�������(!�_�BX���������n�K�Y�y�t2o/lD���l�l[��SR����퇫�EI
rRĪq�dQZa0�SSq����Z�;<XK�ha�9d^��5��ƙ4�	���� Afdgaz�,YӅT�����dM�QQ(:p]�bM,K&9�/F��<ܽ��o�aG|�y�z�Ǎ��fbJN���mۆM�6[��=u
M�-�����u ��i���iBPp%N��I#<����7^}�>�P��^HB(������=�P0W�jw���G���0g��N
�UL{�	�����ാs&���6��d塺@Y���:|t����Š�!�E����)QX4o�ģS�Nᥗ^b�H����s|5�`��
�u�'H�3���%2��x!����=��)S� �<����`��F�u��s�a@8�'�����>�'6,(�C�I���IS'K��+X�J�H۬V�\32�
$���<AC~ۋd���q;�|��K��c�	|7�p�fcav�QL�B};�,Y�6�-���pk5h�6�bs�����(�m��RJ�0�,�&�<��M[(����u�`�,C���f�x1��^{}}}$�-��ř��ȝn�:���!�ޡШ��{Y�V���B��OwJLe��Ĉ�����3SQ�I�0À���ɈFf��{׮]�Y[8�O�1]bSvO+�&8�%��vv��7�L>�4-��$��T,�����g���Ѽ6��P޲���֓� ���LEc��fsbDPf+9R�$����Ҙ���51|o߀e�^!I:̜�-��4~�Ν�r)S��|!*~ː�@8]kHl!�TС$r��x�?b\$&Q��x�����vYI�����{��c�Q}���B�<2����l��ux|�NԖՊ���\��`�X�� �W�J@#Ka��Қ3o.N/����~]]�$Ry�iH
/BC����$^�)J���tW94'���G�+Z׬�����?���az�������n��p�.X��;�e����jQ���Z	�LKANB�֛I�J l�Q:%rғ��B�؟2�<A~�
[�m�B�g���_�j����3y���db$��u��=zT ���AV\��p�5��C�ʃ܌DZ_ �/��R\1��#צ䎥�u1��3� �:>�aוH�My�S�$�˗/��w���}>�bB4�����\��:O��:�؂�'Iʔ��-�27���ޞ^�EF�ű��H21���Zy?+ ��MYc�WjpHP"5!F��K�O�<)w`e.���\�^��5)\^���K�Gme����Sl���'FQ���k��R�@}ȣ��U\	�I����Sc�p�e�����5(�
����v��V�K<A.Nr�NK~;n\���Tx�еJD���ߜk��b�j��Q��� W
�m���?}����}��a �{�A�/TK=����%�`���ݗ��QA���6��5�`.E(����X	t�@J��[׉����!-�r�w�}�af5�!����u��Ā��:8V���rrhw�`YBۆ�����-�@��O�Juق��:���pY��D����|_�0z� p9}�Kz��{����0 V
B,,h�����5ea-%��;i�<h|��XK�W�9�:����؛�{����8씧8�\���������/!��'��i�)��}���X9q1��N�P_�jw�)��Ff�qXOLL���o0צ���M�R��C��;)	�Sk~'�D�tW��p|%��D����c6L}�UV�v��a�U�*�4�r��^�N�db�M.ޚ-�=Oo�	z>��D��ϻMNt�(�NEzz:"�]q,��%ם8��=�)����b�F��Q¦PKi�=�շ����p�qM�,\��O6�=h�����ڒ(q�0V�F~���+>�
	̸��� ��2q����;?��w�."8��}p�)��B��Yݨi�cf�4����P6�EEF���q��#�&�G�'�����)��mX`���K��]�b���={�\�Mϭ�0�J��݃�is)P~�+Ic�����L���66 ��U��O%�����
�`W�J����A��FC*�{x����%��l�����cٲeؿ��.q.\ ~����,#-3�Cp�|��٘��.�x�:�a�:�;l�-s� ;;��@Em#�\���"�c�� &6Nji����F�]u8y	�q|��[Ɍ�uaP���rD��$���5��g���Ȁ�hjmC��$uAëf����Pd�p����E*��z=v~�V�^��d)D�R3ӥc&�+Ŷ��S���N>��gS���r
g����K��j1c��Z��\Y<�&V�6���:,��EAA�Ν+JȊT^r
�/
���J�Z��ű�<W9X�آ��J��bs��Sb�L�V�^����1v��
mnz�Y�E��6�����Id��3�>� ~��_I�ݻ{�⑛7��Cu����}Z#�`4�IBg�Х�D����<!+e��Ipsб`��N���{�;G5�.u\l�$nڦ�����;3O�G��?���Ue����c�C�x).(�P�������ix,�_�B+[���>�2��6l/��-QC���C��6��wO#3+w�y����U�-��$�͞�#����W��9Fh�>6�4�Y��Ox���C�슷�<���B���Al�u�F�9E�1�s=�� V�E�z��'۱�D��?Gv��{��K�PY�I!.ܐ��s"t.~��G^/ˢ��hnh����~&ۣ�7>���hTg��(��M��N6l;���(�췿���5������o���� �����~�Q�P=�'�A���ȧ)~�q�z֬Y"ރG����U4g��gh���k��i�F������T7wK�W��C���h7+�����JCTL,�|�I���ٳG@9q�X����dS��!~|p:QT���&���>�(n��f�7����]�{U���O� ��=Ԅ�̃X{�R��*6皚i��۵ՕU�6#_�V���=C�Tu�:�(^�46����@��׿���.�����K���::v�ă�CT��6�GZ�	Q����'���'�s��[��C� k�	ύ[�g��rf|�?�{�R���?����,�RGk�loGVN��Wt�[T@�(���O���N6=�e0�������\<����l�C��<��[������,B\T8
��A^^�~�mq/���İ�(���>��01��p�0P�����8@ԸG,�����yO[�ڵk��v=^ܰ���"�Q�F��I��w
{,r���zS'QgàPU7�E�E�D�t��}=s/2T�%��9<\�4�����<��|V��ؽX�l)�������f�͛7����?�*O�b%u�Q�E����k��$����o�y��`��!�¥eЄ�l܁��]R�:{��e�u��y����4�ysfc�ĉX�n� ��[o�����4�Y1BQFm��I�֬Y�'�xBr�yԞ_�16��WFvC\�	"vc���[G��99�������ơ��$J %%�|�ь� -��c��/�)��{_ɽ7^����b)LO�Cp��˙<����ԐG�[��pn�.�c�op��u?�+;��R��A�%��_�T�O��9�6�K
%���?�Nז-[�^__/%��2È�[/��-K���1�PQQ����������B�������;��/��~�_����za�!.2f��p�NO�����X	yK��y�K���ݶ�Z��p�s�=���k����QUU%���lο^�e����[n�E�8qŃ�b�{}�gX��	6������l�A�����QZ���+"%5E��2[`Z����R<�dq��� צ�<����38�I�~v(�+[�q���ۊ:ƻ���Ĩ0vj�x^;opX<=Av��� ��w�fwbRJ�����A��]a,���a��M�J�U�g6�@9=��51ib��0�w�}����K����if%c�c�p	�����j���'��������_���a@������_5�l��48�x���+����9�v�t$%&H �5�_$���|�� ��t�xi%���>/�ɥ�(z[�ԉ)�@	[��9��e��_Cy��ٽ���k �}/r)��˚?Nb̠��[�җ������݂�da�5��?$#<<LX!���-eT]�<��4�ʚz|��m�~з�y�9��^8�zd�λ��b�hQ!8�a��`��|/=�X�D�{%��]�ES1wj2SE����el#�V}'J���T3�6a�+d��X��c�E�/˛�*\�m%Ƽ�dG��J�|qEjE�r�d���dF�]�p��ε���PX9�����wV���X89��i������Hى��N�fqb�lFGW�j�e7塚��<�Ϯ<��c�u�J�@g���>���|7?����#!2hgC����R<�X]�(Px��0<���r���F\�I�:y8o�d����g���`���@�����[�NKV#9�E��`�-=�PJ��`j��A%v�:�r<�	� .�W<�8�M\���fŹ1>�Lא�����o�i��&��A��V��e��w�8�#tDE��0�[o���n�[j��x��Mf�iSR���-�NLJ���k��yǩ�>:� uTh �Z4���`Ɗ���<K�y��w�ԩ��D����~��a㲒��v��>3M|P�r�eu e�
�����H*q��Eh������]]������J5���Պ�+gG��Iy#=6 �fD�q?]�U	8F�ێ���]|%YV*&�����h����[���/?����K�&N�uw,�ؿ|IMs�|�����������j��AZM�[[v{fg���{7��o �H�_��,�T(��v����C�!\��\�s�s,a0�w��3x�3�Yj�(R~�C��/������"|H;[��7����gz�� 3;X�_��܇c#?i��~�����m�o����H+I�3�B�:m"�v����T+�7�"W��T�Y�(��}��A2��6#5bQ���+�g�صٝ�-mM��]��ܜ�����`���5��&���ge��>����-eM=A��4{�+�D���9{&��Ӷ�4J��:<^���N;~��YAnS�pzݬ��%>�ʀ�NE�t���*��m�C�V���xlN�W��f����֣�)�u=1##�a
A[�N�?q�&�+f�5��A�/��z=Qĸ�o~c���m�OuSN��F�w˺"˟c�U����������[�m�[�Z��
u��m}�0�@�b�k_Y��)5d8y�Փ�w�=/�s��~l�R��dl$��q7�G�����M��/�&D�vI�T���Q��؊�E��	
E��A�۫�X���w2�f��3m����h$P��� H�4��e�+K�.yF�sq�6�i���kv��q5���qa�e�;m�>zW����/3tJ����UM�Uc��s����+�A�fqZ ���tKcZ� 5 |���MF���P���__�%��q��ߎK�r��o��Ʒ�\e�[@�����lS��?�    IEND�B`�PK   �e�Xi�={L  V  /   images/938ff297-106d-4ecd-b830-d3af457c8fe3.pnguXeP@��B�[q	�ŽXV����E�]�{!hq(�-N��"ŋ�~���f��ܽ3{�Ǚ3g�ZJx�T�   OE��/[��r ��;~�_�+y t}�	4�L��!���������������弄�������K7O���WT  �
T�������z�E�wO]T=ѹD.c��������J}����3m$'ߣt��9Gp��"��ՃX8�JDp#��Mf��\(Y��s}g��?�?Ƚ{x�����F��N,9��W��S����ӯ���`[*91�=Bq|
ܛ@���^g����ñ�`,�i����?�v��w���%��332&��b�ζ�`J999����48�X"y��t�����������q���y���/.7��{�g�7z`�Ư�И���CC2�BT�a���mn���ـN�?�ۻ���q��ӧO�9-$߾}��+�hhh��T~������H/S��k�aPo*��]��+���QXX8tpX���qr.�H���`��C���XM��'
ϯҭ�>�V��99:�)%ө%і��)��h ف�s䍷:P��Y�������^��www�A�p,���%���%�a�	�*�njX���-Ah�d8�����ҵƘ~����%\a�PL�R�a
.lAOۅ�k)N�!R�$�`��,H���PN�cc,&!�����( ��Xa\ɾ�5+���M��(�%�K�7�H# z���ѰH��QZ>���8��Z�T����?�\�WDr{ދ��|�6��z��9��
%	�WHP�,�R;��))U/..��Y��#BdD��鬧���R�ɼ��3h<q� ��B~���VUU�}���(��&� z�1rqq8m9J?FTTT0�n]^\��˂���T���[[[#��z����6y�t���,Z��gB�|���?f*m�=�������W�I����,�R9X��Р�j 
�R(D����z���"V/Yp@7�؛���	��3tg��YYd	ʫ�<W;��nX����E�_���Y�Ј��XÀ-������X��!�|s"�:���U�|f�1`�YsM�j�`�b)�*�-(�m��@-�X����5}�V*���:�Xz7�"lA��{~vV�ʪl����sJ ]6�Ex�.>"Ü~y)�LV݇׬��<����x���N�v7���9�zn��N.�h����@�!ƨ�u%���RUK�����H�$��3D[��e�-��x��Bm
���m�-WX�v�����-�L���<���b�¼�?��<Y�[�����2����o�gg+�G�W�O���K�v��zWC�\.�mC��xڑdB���gG��H���o"���s[�xoٷ`۱,劉k.q����,n'�/,�d�ƛq��e+��ᄶ�B�t�M_���4�߲�s��o>��\V��ű~��*��]��U{�T$9)G:��>��(!d@���������N�kk4>v�
�oZ-O.�p�g(3�/�~���v�YF�4(Ֆ���qY���.!s{Ę���4��g�hȿZ�Ӽw�ѫ�� �V�2�|�?�����j��䉉���Z����$7(�5aD�XsOYۧ����)�X��s�a����ddi2�R�(��b	g���k�fJ!\r|�$���e�C��$��E/kH�[K��D/��D_��¢��u\X.k~:�Tx�՚bߊ���QDC�	WzN�l#�rQ'樓^&%S�:�(��e(�$j�5�q���19����$��`0z~	KZ�$��ozc�~�����osX1+O��Ac*!��}�򡀓��N@r����2�z�)��u̟Z�;x>��9�}q��� $+�L��+9��B�f ���v������x��4�{�b�^�!���%�8��|>�~�{�`�ꪗ�^�U���bX
���Jf���ATGi+Ț������ 8n��avC�ZF^��`)bS�C��+��!���w%ֻxt)Z*)�$SF����x�}��eUr/o_���r+�*ٝ$f�+O2�7�(Zd�'A��pR"233���M���8!zz��9��yP7�_�_�����0b�̥̒�ݴ��jK��8<�ħ�t���F���D_��A�8Z�������'s������m�%�Z8���$pvZ�ܴT��6�N�}�\�M�Y\V�_�k`�,��Q� ����k�
��w��A*�g�R9��NG�u�8��9Ƞ2��/
t ��3�'��I�l:��
[��n�e/�OO)�w�GQ��r��'��:�G��S&Dm��z�݊Fѓ���p�Ro��b��Z5�db�` b5(
,���a�ǑI9v�%?�B������x-�޽`���Q�,�Q�C��t�2��Kj�1�?��#s|">�����'��S_���u�?�%4G��C'��/E�����@�� Ħd�1�B1)`q	�����(���c��\2nhPB����aN�YR4|���r"B=+HC+�����,c `������=�&�?f�Wd܆ş����7-d�S)���$�E�«h�ʕh�|�`l:��R��l�P�K��f�+�3�B��m�,�Qgт}�ݿ�#z-r�H��(y�eb�2c����C���I�$fv{1�����=��F�^6�_��-	������2���Y�k��OhN���6rc�f8�Pt���j���}��pRCŽl�`����E2�9��1�?QS�@G�d	�}��ⓞ
o)��1A���TY�{B�]�y��� Q{��o�mMY0!zR|n��mɨ(i?�t�Ui[�����[yf�$Y㘰u����Y�B��!5��75�-��#�w�YLc"�|�G��ΐ,�wwWqk��F#s�#�wە&{I�le����V�h�ŝ���(���+3�Hlg���:k�Nxn��IT�a/,�pj��ɀv@��t�qğ�~��B��L@YVh��=F���s�upߌ��2�^���*��t�N--��s(�.�58!�F��'�r�?d3�{?��-d����-�r���l4��E��h��~/֗� �{�c5��J�wsE!��U�ͧ�,��hrM����z�h9���H�C������Ѓ�zXmI�n�!�2�c�i��D��D
a�N�6	�<߀,���>��N���k�'f������Y�Q*����2�����vdr�+1�K�Ⱦ�Ï=os��S|QK��5�)�$�R���|�y�A��"�
��Hhݻ5pf��Pܭ��,�bJ����`�4R�w<��g5b:Oҝ�<I�,whS� T`�כVarz�m���!Ś[�e����m�e ��|���'sI�Bx`��,u�]*\MX���^J�?k����K��w���) &�
���)�´R�p�f�]T|�z$�촽��2@~�K���s�Hi�L0����
�7`@5���	)��(�k�{j�Mb=�,��ߜ����52B}BE��c>x6�DOkh�0%
ɖ$B��U���H^!��<6�>���KDs���u�&c@N�#�lĞ��ܦnƉ����7p����*e<)ѕR�����S^R���\�J�[N�N�(���7Z�%6,�Nk>��ѵ@qM?>4eQ�3���(ӣ��1bp�����e�,�QK��𑐁B�n�2 �'�/������u��.SƢ5���8�0j��IJ*�t'����0�-^��"E&&�f��2{�~
o�%���'�OY~����QVb�UÉ#�Bh4F�À�б�e�D��L!���0h�A@�E����Uq�,�:e�(ľ�zc��:ӽG(����,�^�'z]
O�Tٗ�bl�}����@ӽ��,S��4g�W�F};L�+���io.5�N�������h~�oW���^ʏ&h{E�ζ�Y�Ob�J���K Ĳ�jz�� _C�]+����'���L��b�����_#m�P�3�)� �O.F��<�="�=+�zf[�����6)�Z�!6Gԭ�	٢�T)D#!�{��	`,W�CWx�7�a�ҨQc���e˱r�҄�d�4��IINhє<}��F�Dӌ˱�fj��}��s��1�"�z�Ϫ�3��5�q�fY|��~4����@��R��e�y>�L�S�N0]��h����威[#��2����MZ:���V�{��I�k���{�OL��U8�i�꿄�v�q1��1�N�ec�����_�g렌I1EH|��϶�זw���%��Co4U$�Ҿt��[�9�߲njjk�����&����Bv��>uw?��`cO���1%soչ���.�=^T��$=��PQx-!�2��X�	S�c�����||l���^}V��{_���!�w�H����Rx>rS-f�T[��Wq�E����Q�j}Tr��nLl��D�p��D��Ww�+��<�9;?/�-fJ�X�:Y��By�s��v�(�}��E\�)�i��ځ�H?�䝊�KVn�_���pD,ј���d��)����[��s<����3�^RϠ�!t��#޲M\���ҁ0
���Ыr3X��Y�-}�z�C��\5�@j��=-v� �'��B�?�3R�������8�P���I�(�ԜF�F������c��*."Yޞ��3��ÿ3�s)L�hĊ	�:e����Cx�Q��5�_�e���Oa�]��^썑�C�����Y���ü����#<��0-�l���p	(����_ri����y��~-]�-LD����G��^�q����[YDo����?�\s��ց�ߧ�C����q��/��z���D2?� E���Up�-�����y�E!��Ty���Q� �v��J�3���	�pJ"eT�1��f�T���@�>�d�:�3W�����gc�C�5�g��!:]8���RH����r���5ה�������Z#�2�$���YJ*Q��,'�Ւ �T֧\W[��ī4W�,ưx��Heu����7Q��^y��=\���+��b(����vX�3�^�b�4"(=r.u&SmmkC
0Z�5�S��D���. �L?���0,���cG�Sc4Xġ�]bT�JK�n��)�v�oS<�GŸ���K�^��7�Z��cUf����)���h��K������X��]�΅�cT�I�� ��}��،�$�O6O(R0�#�^�q�r�s6\��]�a 8ᢑ�ɯw��N/��\�9��h�]�xK��2�?�ْm|�|ӑ��O�A)�{���g�+4ﾟ�du��V�1gZq�BZM[�i��3�S�l�PP��~�yC6'�Bk!���~͢��T)��6#/SN�kg6)Y�����Tu��q~��y��xl���LΦ�}��Y�����_!���ὖ�<jν���G�� L"��Uȴ���#<�d���˞���Lm+��������b���yqp�SV�^���͍!�5:�ds�z�����[v&4��_���VE.��j��$�n������Mi�.���I�IG[�銾�P�	i���=Ky�V/UN
Y����zc�������t�E���%�������s��ږ�Y��q2���fǪ��wf����l^�6E|�<&��{�.=�^�8�"ѡ� �q����3�xf�>�������5Ǒ������4&��4�!�}��*e��Ē=rdFd��8�b��z�P�n:����p�x���v [�u�ׁ`�y(� �T8H��4�f���:,��R~��y�2w��,��tG΍��=��'IR_�[z��(�Ǳ����#b��~�+2xW!�ƕ�fIgC��]6�mZ:�j��6sͽ���[2��GǺ����I���mf߰r=!�ĵ�"T7@������Ռ&b��[���C����!�M��m��#>;ڟ��F����KnIzYu��[Bq�xA)j"�0��m��R� S�/I��G;6��/L�m�Ы�X����B������ؑ�o����LK�����I]�j��a�y��`�� o���������+�f��O��H���bphV�߬*Kg����]���*�C�Ú���}�u=q�mE9���"��+�`g���D1������mqu�փΎ_���vr�m�q�^Q�,*�ӷiCLC�x��d��]?ه9�+�Q!P���Eɪ*��w�K#8t�9n��x�1�jo�݋PJ�S7�Z�X&2a���(�p4�1~�����fh=��g��:�b���p��H`^l�qv^�SO�^;P�C�������cA�c�U�k�G�|йjP��C�%�ѯ��|����s��M�Y���8���u����g���-���&M�
nn�n��9���`�����b�3dW�O���&�WɃ�D��ݠ�z��H
�����T�����AىC� OZ�x�<��LV	Z���a���A]����zF���t&��7�
�#�����Y;�ݬ)��9�R����P��/�=���wl���b�խ�GJf��F\+��9պ���Q��J��s�0.}����E�YB]I�{�U���މϋ���Z)ʯ_W���)�Cu!�ƌ�1}��}�I������G�an��'��|�Uη�/��/��-e����W�t7�Bn��
s�魩D4K&&8Iٍe��W��=Ӯ���/i�[�^=ܯ�ji�e�+���ե�k✿��z5�v9���?��9�x7y��� =�7`������m���d`@�k&�lii��T�2\��}���@��;D(z�k+�.���Q�z��U��X@���L�Fr����=v!k����\ڀ���+���k��Z��=�|����N�:�9��9H<	�䎥��m�]C�V��
�𕦧�n��<d��`*��4��0c㳴�M��L�������c:&��ˢ�����t�׭9���c4 �����R���Ǐ�byy8xeJ�e%!��D&yjD����.8�jV����47t���!�!!�6fX�pQՐ~R��q��	��4��-�c��T	-���[8{{�k׫#r�Mr��#��E 30XM~�������[��|ӻ��-K��yhnf�d��|�g�g}mZ��%R r��%Z44�l��+v0a����zn��0R[��n�}KEEF}~>��w9�a`O��f"�7�X�fE�Lv���q���o��z���c'�����"q{V�EZ�D/��t�xD��g��E�6w|{#�9@D�M\�:B [GP7�e����f7����������K^S d��J�"ܞ�;xI��'��"��&��l�)8@����$i���l�gJ��D����XP�ʔ�M6FA<׷o
�p�Zca�S	��@.��ͶI�����G+G���O�Q�ռ�{��7��ד��h%	���:}0�RA�侣n�g��ו������I��%k�_�����s�Y�����|��3�@���"��WPS�׃��z�|߫��1�#�>_}����뮡��ݒ��5���7'K��H)���=E�_��Y�����]��7�\��H]ݗ�X��Z��E�<�#��"ě�z{XSsG����=Rs�L$�=������_��*-w.0"������D&����G���Ǹ�l�'��H2�=���;A�_���q�eF���e��6��7�[�n��y�R��D�Mؓy�|��T4�����PK   ;j�X�&�}[  y`  /   images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.png��W���x��,@���$$��[pw'h� xpww����]w���{��p�sf�L�tWwu�S�]���(�P@ ����2s��{����[�<�[��)Z���@tq&����醌����Q�ܕ�ã����0��Ќ�P"��b``�E��X����t��a9�檗�����EV�����*f7M�?!��ģ��JHH�`�s��m+�>=,?��8�B�ybѣo�h�I����7�.5.��}7�O�3�����1�]��fPz���	l5\B�zB���Ǡ�9�WQ���t��ԇ�t�D���=$9���y?����K=�`�?y.��d�bh�h�� ��;|4��e44Z7���A!Ɂ��Lс3N���R����BS����d�����_^��Fe�v�����t<����)^�"��y��(�N�Eİ �7�R���h@��`�(
��@�� Ё!ğ8��(	/�e$�A�]wb���?d)-g���#���(Dr�����C�G���!I�_��������{'{sK��.�f���P��z�>�7�Pz/x}�^�ʧ����f+%O)%�.V�>�9y 8�o�Y�ڢ�d4q}�o����V��؂g`�`࿘��u����_*�/M�ܛ�C�M��T��0=��������,�.^��_�������8&3E���1]����ߤaV*宣�K�W����?��P��|����������gi�j��fJeSk�$uQ��h�/ڳǠ��S���+M�x��}BM�9�+��rE�4dMӌ�����b�hp@���/fg�����Njy�|W"D��=P� �LC��˟@2b��+�U��=L;S[�1}?�	�c�'�z�ײn��Q��I�g���)�GD�!����3KWEc��Ǝ�YXG����w�W���qO�t���?�z,�����=#�Mp�����9Iq�����]fn�����\QQ8қU��X-�?�瞭���ܷ�Y�}x0���]���Y�c�����MY�W��Q����G�E\ж�aL��f�y(�3�_������ţ����6����)A�X�֕z�ΉJ+a��©�����\l���f:-��¹�/t ���'"�vy5��S��Y��u�èh�z��x�ۣ�ni{0xq�ʇ�|��_#[���%����*��5� ѬXX�'����K0y &�>�NTm��Q�׋E��j�@�	�����z�f7�*�������i�ǐ��	z�M��)+.���"}Ƙ�s��̥�b���93�R�R /�y5R��w�>�v������Fdt���v8���ډJ$J�ݜ��t�+�~�?<��la��綖Kц���x��+��0Z;H�fp�;����7.�c�sϋ����?L4j�ctҲՊB�뚚�&�n~��/H�X�A�uM�Y�����5�W���a奫�r��E��泑�'�'CR���:N^��#7�2�d&�o�ȩʓ��_���ne������;]V�	�%�R=r�G%N�UH	�|:��}�$�$SX9\:�H\�.)ah*-Ywkݸ��l7��TrCnElN9�����
��xwy�����=����$�a�V2?�I���)��5V��'<<'EI�I���%���-cO3:�u*b҈�Kl9�@V[�~%M���0`r�b$a�k�G�V����;-����m�'�{����6H��ca)��rw�p]�s'%���R�զ�ţ�L�L��Iծ���_�me$-:���y�'N|�ޔ /�B����(������\���y�I�f�f�~�ٸ�(ka��o�e�����{�)T�,K}!Q��`@6p���5A�`�҇��P_�3/A��8yZ,,,.1FF�Б}��'?�-_arFF��#��k\����~y�STf(JKI��efe�zQ<o��F8���>�!�lU�{�)�p�w���,.vj|?�!܉)_�1���ϼ��+{HQ�W�gmq��@WB�`aVN�)A,��<�:�^�Y��CJ,޸��o(ǜ ů��gwm�@���8Xt:U�.�3/_V�X@Bs���8�&�3�`^?�k�of�Z�0���%��2IL�P�������d�*�5�-M=���m�D��I@�)4�
�wQv".#(t"���k���R��,�WR�	 �ϓGEe%P=|��^;��_I+[kRk����J~��(�:I ����|8��d��%���z2=1�+�u���k!�p�P/>�/#�e�4�������5��D��t��*ɟ���8L�WD0�OD�(ɀ�6�a]V*�,_�r�קbC4�\ $�1�xJ,SR�r��z���oTgdS�[���C���m�:-���5�t��I
�KͿBʜ^%�*��'�����4f���Q(`���u
hR\.
���쳜��dMV�#�������IW=��x��1�ʐ�ߢ��3�����B�%L�D��!4�0+M��f�3���o��&x��-����Tl��d2��%E��`W걆���	�ε�O}�!9b��7���ʷ5���$˛j.�����K�8�j����#�psJ�{"��<|��[�v̆[�mIR+�?v��psL"��kDs�X��ݕ���)����2�_0E���c�3��Ȫ���ϧ����t;�	
�UUUlbb���n�F
66,�jA���IL]N���ē�E���((s�ak,)d o�~��oR��}�Ku=<��1��Y��t����K;y�V"(���n>��0��W+���,�P���sB.+ܚv�iND7J�M����w�r3����'{
���k�����-���4�j�cm\|\Ѿ�o�s(��+�cz;�7�������ⶳGԡ�5̙�~����@8�.c��m�� XE]m��� �0��a>�7}eY�՛ł'�äa�.<�L��ۄNm}.���0s������O�TUL��#�\�������.'z�	�:ڽa����H���x:N���w�ng�4���$�S����',x@���2m�]ەt�QO�ϧ��zkZ������ HS�f���`�eg_�;��l&F�� ��۪�� 0�A~�����{8ܙ%I�[��������灚��|��<��':�N��o��P�4L�Q�z�������4�c.�{6�?�2 ��U�Tv_�&y��v�G	?����W���4�apP;A��U�4�K$�ԧBG7�%[��r�6k�n4l4��i����=���d�0�����V���`���C��s)I�=�%/�4�u�9H���Q����'�,W��ЮY�B^ī܀��;��@��T烌(�7���v���98��Zݾ��1�����78HEC�xR�����J��	E'��=����Ϫ@*�^/+�:*��-�C������r�(�*�~3鄖>{�q�/���f�H�ܐyV]/�����ްd7��r�ߦ��0 �jfjn<:_���2CYV��Ç]V�v��+t��%s��k
/�w�{&[�s\4�)A�k�=�v���-7�#7DW�������"��yZ �2n����Ir_�ʗC��62B�̘�<�t~_�����Q�l$Ȏ����%>�=v��TpZDD���M�Y-�IF�/�pq�{Y���<���s�OW��Ef��iΉN���ߥH�:�0���(�8�n�5;�����;w�+�O�e:OG����\{�B��S��h8B�ޅK��NC?:=\K�{�����x�?#U9l|^}��r��'��c��)�=�Y��F"�쩅��h�n�x�ﱿ���ܼ��B��˧�pPx�����C�!��Gx��|�%���5Uq���pH��}*��^�{V��cq៞=����U>9��e�~�	��b�u2�++��pR�ȼ�굺�9J�ޞZdn��w��g�C����R�sB�x)�vb��/WS�֘Em?`�r,���]�<��C��H%�>�b��)�13tɰt�?}�2���x��iz��V;R}�s���7���&g?)�]�>^�>����c�����X6������I~�I�%���5EA�N���l�b���ͪ�\�N+>kr� 77���H=!��<���,�-0ߕ��D��II���"aK[|�|�3�e�_��z�;�hO���a[~���`�Lb��e6#H����M�M���*Hd��.^�$`�8�{=�r�w��K�~�y�b�x��>o\>l�{m�`/�y-w)�z)�ym����8I��N����[ �:x/�=<Ui~��.��*gM�E�77��El?x��{�&&nظ`X�iؠi��n_ن�8�p���n�t�Ab��K�Pd\;����.��o���BU� Y�%F��Bp&>�ß���]����k�k����ֵ�}�APy����5���K�M�K��k���r��jIy(C��EO��N�/��+��sU���ؔ�¸������Z�x�<A��u����d��:����t�`����zC�W��_e�.���������vY�S23cA�r����(hi�ظu��뒦/�T�չ�Z�M?ub�F�(n�f�-�u��>��f'L�������0��:����d����!�J"F����g��ɜǒ��9�*�a�2�F���������d||��>��hd����T��cw��J?~\�ή�Y��no�j2���dd`�n�>R~mH��D�ݦo�>?0�#�����c��E�jR��� X��<xkpE�fd��
��b=*�2 a�SW'@#��E�������|m��R~L.D��8��\��ݿ�Zj����'����ic�����'�B�5�% ����0���[�΅ʒ��Җ�3�I�R�R�_����)8��LLK�\����o�!�����~���x���C���?	E#z~��*�f�.ɫÕO*�q��ɡ�]4�+)j�n	�ܪ;/������g1e�I��Ӣ	@����n���v���}f!S��G,��"�\V�[��X�|
fa��"�L#K(i�X���|��S���r���^������G��R(���O���moMR��t�Z�8n>����U�!¯﹣�v7��76I���x�y_�B�������n���>?��|	J�+č��YSF!��8�|(��|f�C�V��d>�{�U�w(�xx�
�ď*�i��=Ճ���,��1B7�}|$������8%�A�G���j?�KȥBIy^���m�7�-.�(���EA3��3Ӭ��ot���m���Ә�N'&�2��ڣ�e~ge�'oY��/%���$t��j:�Y3ꉠ}�F��殺!��`��xg����ua6���T���w��j�2��KX�Rh8��2Yn�F�Ie8y��2_�&/))�R]�N,��M� *�� ���v{68?i=5�nD�2��ed�:�'3�h#"ƻpz�Bと}�R!&�����'4��[�oڮMJ�����������b��$?�_X�78���؋�U�D*�H$ǁ���I_�Dz�ɳ������]\\�L�z�����̒,eL�s���ꏈ�^K�G�L�?��.��a����贼�6��z�"��\�ęq^�_�*��q�h��{�c{����y�
q/mw���0��2w*�`��Ĕ�/ Q�4�����;M[
��L!X���kt��k��
�,	������D�qh�?4���r1�U<��֘썫�M��d�q`�+o�����4�3'^��S��$�vUGGG&9���Ե�`����_B`�����
�V��@C=��d@A�mk=�:i�ޙ���A%�oe���^�c��~_T}q$�B���".�g�de{��qX���.�􎏅{(~�<����r��ŢǴ�?L	��7��C�fo/,c��R���&kπw�o�ӿM[P߾Ϥ/���宥34N#�Me�O����l���O�MFe��z�Aڊ�G���p\H$��g ��4��[&�D���5)=�gRS3��}�
�f�fn�V�����T������bꞘX�.�g���^�����$2G;���M���
��`JJj3����2{QeU?�rS���fL�Z\�����tfV5��	�wk
"s�I��Ѳ#n2�_S&c;?0��{�6�}(��r�KZ���H�|;��& �����kdw�6��>�tC��-Kwк��R��˵���v�VzWhi�џ$^҉�	�:��l�s��am�ߞ��Cn4�	!�J]�����X�'Zī_��>�a�����zQª¸9�����B/n�Y^��.>��������4��� JBq���P9�W��+���'$�J�Z�T�L=�J�2B��B�x[7��_��/v�aTv~�K|闦k�g2��W���Z���صh�T�{m���:ָ=�/��W�%x�dP#G�d��(��4�K[�%���}�W�Tg.��� ��|<m�����P����"�y�9BIy1�s�g�Hv�v];,��n[���D��7X���?vi3��b��A����>_��9�ȸP�#�:8ty������/�+:�g^�~e'k�ħ"v���Z�����Z��{j�#���_���
�d�wJ�Q���N;�F*��*`S�"&��V����{�y��V�Hs�y�b�8\��~/7V���o*�֎j6v#g�{�#,�E�,��-��d�K7
�8nFA(�k�]%��TA������	����E�ʭ���Z��ʦi�D}/df��vB0RǮa�qw.�rx�pZݹbp`��<�Xx���I@�"W���b0;}�n��ZA䅤q���fM���~"onb�p�K���a��#����V�Ksj��l�Y�W�cBw���!ʋ6�\���3[��������|�}�ƃ[+)zP��,�UC�R�?9ϲ��=�g9�Rμ�|���@B>'ܚ�������EM��У���*���Gk��-�U��7��MwiF�K�����*,��ka` p\��;ط#n3�^�̗����D3/�%'�e����&�*�&�v=TWm��`���<_f�����֣L���fH*]u�%���tj��ҨԗRP����e&p;��p=A+V�2z�&��56���cf&xI��C�%?c�A�<N3�7�ԸEHij�R +��@s�)(`����,q.lؚ�E�*�۠��[����A@�����s;Rh ����d�x�g-mup��o��h�N8󜳿e-��~�pvlv�JL��aI�~��+aӿ(	3O�I�!3�,Q����#Qp1�;VW;4��}�(��O�Ϭ�z�/�,/O�|�i��%,���h��ƐF��>N��@8�C� �@+* #�\ ��sz�%����Ca?�����]���Ȫl�0�
M6�P��uϐRn�e�A'�W��B����څ�U� >�,䝚ʕ�=�	P�yO(h:?�]�\�@��zb����Se@Iy�y��yh%��SR���_:I=�(kl�Q���\8Ԅ~^�g씈�Q�v��_����AeL ���i|��d�c��ijfƣ"��/b���j�������(���{��q���Vl����FiG�&!��{��s���en�Տ)T���hZ;f�Z���ӵ�w��
	3�"*��l���22��)̫S�gѣi\s,��vAM��U#�r+r�,cT[e5�5��"��&����js)��ǓQk�Ro���h�6�>d�{d��T9�b�˒uڔ�1[���Qr��y�t|��e�3�5��l.����kA�޷{A�}W��}m7��}�;_�î�1PcE��.�k\0��Z�	+'h[�'��"w��O�^��3�#b&�t֗�Ǆ;&�*�H��'�]���i������K�C����umm'M �\�M�3.�%�G��2XΑ������H虙�d;`�[�Gq+�п'B�fk�p ,[�u��~PU�ɩ�ڍTc���eq�ys��9=n@����`�S� ��-ڎ͞�s|��9�)o�` 3X������ܺnG���;��RJ���ݧ��8���[;���+t�[�SR��)�������%w���ݜ,�=��@�����3�j���-�x��6�.8��4ᤎ%,�4f�=��30[�	�g*<?�����ɱ���UDw�Ɔ龠f��Rѹ!�Pg&�hg�����xFg���V75"�Y>�->���Ѧ\�ݑp�\�������Et�R�h"���:���3E�͑�ne��c�g���4�Au���˼,��-zc��429��/1"FA>���JX�����iX�n�]��g�����E�I�w����#"�?�yYY���t�H��u�K���sz@J����=�{Mm%~���lg��I��5݆�%Ɗ�0�3��FcI��1�`Y����Z����2��b��y'~;G�4I��[��eU������׎Z�G�*V\e�zM�s����^�!T�Y?��c����_q_���Z�) ��村���!?���w<���S��t��G�9�rc0s�$�5a�彐��|̯���?�vC������m�<��6v(��ZҐ�:��~K�����>�i�+�Ҿ"E!�$��Q��A���r�|����Ö��:��7��K�����Ճ�P�eWa?׽�u���Sޜ���bL����I�ZUL�y����\��e�۹�"�p��`���x�l�'�K�}!���Na�� x��Sn׋j����BQa�y��V��1_tbn;�A�l��z�����T�zM��0����¾^�2��B/M�8��7��f���n�h�m�tC��c:�L�.��͒��5�',���/w��}���%́�����MO�Kl&�œڬ� ���s���K��\Ee� �������+�k�RU1�A}y��~��M�O��:.h֡^l�!�����[���s}��/�Znv�vWܐ>�Z&{��.����)m�!���_��:�S+j���>���f*ii-<V�(Z�L>n$u�h`��5�A�GD1s�����z5�o��!C�����n��7'+�D0�\č�~�����$"tkpE���:�l��#e�w�p�is?��i(��a�?��8�%$З�%n���"�ܔ��Š�\Re&��Bj2�?���['2�\z��o_������P��t�}���#0�m����J}�"�_���c*ӦF���s�t�ڎ�=�.Ǳq1��KM`��j'��9�"��]E�J�迬��a���3[�ˆ���%�U8��|.B�
j�F폼�e��zk�(;����쪢"=e��BK�F�k)�������_	\c���B3�/·�bM�x��5mo{�_�b��KK�$��\�zHaT��& �P���9����Y�@�kZEE�	CT]?����u� �c"����������I�#`�U�Gd�R:םqm�z*�(��H��QaM�ڮ��2�r� �I>��;\����aGo��cf�d������l��t�k����!m�]3@���mM?U�DH��BF� 	7�wqOD���@�:�w1?��g<��;��%�㚰/�)D�*�#RI_�Fq�?lQN��T���,F�p%A�.l�
�~^á��j���gɵ_�q>���b�%8؝���@,*�H�
W���]]b�����3���Z�	=EK�"��9xk����ۖ�����r?�AYI	K]�3�g5W�F��Z�ZZ��gypE#��(!��=}(���gX~��&�/_�.)�N;ol�ޖ�رk9<��Q��4���N�	��Z���t>5��|�m�W�b!�`.g=3V
���3�z�c�_۽͈K�Zbw��2h�u�4�P��,�V�m��h����t�+]Б�K���� ��T3�|�_��������ݞ�> �$��3qm��-�p�~ 0���E8m%&/�C/4�uM�g��5ب7��=�ưZ�g\�Q��iV�٢E�im1
��NN_�}{��!��t�gy��j[5����v�E�X�ڲ���#��LH�*�zw�Iҕ����������$\�h�5Pn֔����%�E�ʢ~q��k�>ߒӠr/�	Cq�x�m�俙t�q>��M.�r���eu��LS�v/A\>j������2X&�����,{0dOy�#�oY��UJJ��-���q�{�F��CۤE�|YB�o����:�g8����������!�Y�>���c޺����_p0�0�B�0�� �H_.q�-��NP�qɾ��c�-��wD
6���.e����m�R"9aa�0�����IP�ԗB�|`�1��(��ZD�v�ߚ*�Z\>u�=ah�kq?]��'��=��&��Ňg�@�>Zح�JEl�,��@KK�*��h2�s�����eU��~�o{��e��ȭ������T��w�����qTjR#�7�$P	�b��{�dLwU��IS�ݵ:K�4{�D�l��?U�K��l���g��A1�a�D�RK�N�369��d��#9g,OΔ55�3�	;�j5�vmPa~����!���e�-�~l5���D �>6�r i��i���wY>y���ɍ�$��4S6�V�3i�&/I~��AT�_o=5�����1s��]����<��\�F;֖�V��ӵ��v��#7Ss����ZͲ����<Q��5XRUc���pRah�����T� ��KVI�]���'Y����U��+--r~�;t�}��' ΐ]ˊּ��f:���vQ�GWpskc�l֑���������h���/��$LH�C=� }a����Vg�⟕";��N�����J�z��UF&;{�DQY7�'���vЪ����YoƎ;%���[/���j�{\>}��¤�y�M`Ż�]<�"��**��03��ʚs �9ɕ����~�����(~��H7�LYƤ�a���G7ɽV>A���-��56U�K�Y�;��O~$�����d��c��y�'��0)�5�������z\jHr2%K���&?Q��wؽ��%�.�cN���~��s�ϐB�¹sPRWW_)�?�C�M-�z�����TGm��^욐�X�aŭc�F�(Z��O}xc�9����7h�Է��(���F�%��{y�����I�3߰��+l��]��Xܰ�+F���)����)`�Q�<hI��������Ia�S(�D6�c}Jl���O�I^�����1e��y�G?\]_��D�Tx�v�ȫ�Vѐq��>�N���C���mv�y��q�-���Y\BteU���^�=�L�{8�h|A����[�W�ݾ1����)H���r�m�NVr>%��Q�Chu�K�'�7�h~ˆ$�I��e���l���SD	I�Zs[Օ��ދDF%U]4=p/���	!yj�T�_��N��X���V5d�;��k2&	=<F��!����e\���>����z�$B�s&yL���P�$d�o"�K��%�-��D�a���p4�����''6�[�(>�W� /����m��7�_@��o V�R��>��Խ�,�2�9obleQEiU>)����qu�"0)�<��hΞ-�Č5N����V�Y�-ɟ��"&qtt,��|=���X�����-,�{1�����N�A�5��I�|���n]ƇD3;|Y��ޤ��Kᵚ-�ӷ�!�[���y��ɡ,s��	$m+QR)���i`K� c�:E�l�yuU�g���s��C:���R�3�=m!�r����ҥ�oS=�H. �N?�����_�%C��.�|u�:t�H����JD[],����r�z}�J��m{\�ޗ����lU,�m�h� �b)
���h�ؒ���L`lB
���W[GS.Δ�vB���m�<�����|v^��w�R�����֮۝��Yb+ ꀭ������*+SAN��Gb���z����f�V�M� v|�����*sj�Ȅ#mLJ�'�_>;/�KH���� ��_��:p�v� �R�xZ��6��Q�kL�f#I�3P�l���3?�qDޞAVJ5&�g�5b�����Bщ�]����c�aׇ�>��G��%���#	��Y���r�S)-kCp?�ra�ЖE�w5!u����C��y�C��|�5��71Ye#��=y��90�]��rk<:6��d�޼�QQQ��0̖Z��D�`�dH ߛ`<�;:򁚺a��H�]�j�W�ym�>zY��~�}$A��%�\�c�tDMj�\�*�oX��2f=V��tcE�ҘW��d�u�LF	,9�Y�@%SP��!ί�� �=��A��QP���[(�v��p|���R�m/��XN�")��`�+KN�j� <O�'�G�?�SSS?�Vh�6�j6#4�-��l7���C����hpQ��L��L����:�#��;�W�<�&x1��������ؘ��b<����3��z�zu�4Xe;n�m�Q�Ҵ�Ԩ����q���g��lN���t������1<����s��v3޵��-r���5�1���U/���D�D�!�,͸<˷��ɳݶF%Uվ.y&ʀoo����_1�ð~[M�����z�6���A��C�J���w7�ᱳ��~I�=���D�����!a���`�X�eP��Ю���z��tp���ſ��m�@��lQ�t��w���tw2���G͍��d{���p�H���5�H_o��uI��������~��qd�g�Z�\��N79�b���?��Qӌ1���ɔj�Z��2/�I�:�B�VE`
#���Ȯ��芰���]����b����Xma�U�گ	��~���e��	s�%�9�=��^�LT���}{5v	@kҾ弘�<K��<d)i�w�Z��~��2�떠�0EE.�k/�<(�Y'���2&1���w���eip8��k~�uz�DЌ����q��6���7�{X�5w��������=�`7+��"�;�K�F�;(�����!�׌�|/O��G��KR����-{�$�A����n/sɬ7 �T}��0S���,�;��h��rhx\x����[4J�D�糀
��R����j��g��k���F|��.�02��M����7���X�!��(˟_!m*������V���[��7����EN��0�}F��ӓ�v�z���vm/S�M�
`é��P����̯G�X�MfU}�苠�0���\�\~y�`k=#H�y��P�\�:��\aL�J��@�~�jȢ�\���^&��I��/ (�E.~���/����g���EU �z��A��\�(o�Ջe�iLo~C�bi�qq���d�f�H�E���Z�_~.U�!	�&���e>�2�@�_ױ�~��t�_au�	.�BE�N_��e�P���ey�;�6���|���8��'�`c�j�v����3�m��\�[e%[v:�D�M�5~8���X��~:�˙�ͦ�ذ��k���ډ��0��J����^�k�{���J{j�>�3w>:�|�9|��]F�ϭSE�'H��Ϥ;18Ȕ���o���X�ҹ�J��j��[�i�1�F�;31?��x��Gj��	qM����> ��v<8ތ:�A�b);��xq���ص/�5_*��>��&�����A�r1����[X4A���SV7ç�-�ȳ�Ê�N��6�������0F�N���'���Y*��*ZOX�F���7��Ⱥ�xV�����XK��xK]�{��z3+�P���{���Иl��Se0������!�� ��h�z��^x��4:�Iؠ�W��F������K��T/]��^��;.�i��}�"�'+�[E�1=UbS���ff�DF����IO�WUW7~y�լ6��͢�/�d��`;�[��Ubu[��]����JF~oII��D��[��w~�}���$~6�a`�������p����Ȃ��TP�3��s6Fntb]it��mѕ+?W'�O�q��d�w#��v�P��fD��5��V���U�jQ��Fb�Awe�����ȉ5��aY���Ԗ�x�\�M���,7Ϸ9���B]�O_�1�I�)������/���)��B-��������q���ME���~~0��D7�U��b ��gs{n_a�0���7u������-�%��t�ѳ��~�Qe��e��Df�aڻ!j��M��t�M�դ�̛!����[SS��XaTc��6�95H�]�E��;
���ȡ��e�����'�W��ĉ�����.�= m6^80G\\x4rbFJX7�Ka��2��?�lB��g�;�����CF2��f6o�l 2��?������O��C��ͷ�,��R�͘%��t>g �9��W%�����-~8����h��Q��Ͼ���_��:����iz\��i�$�)+X�-9y؉��z!��E�jV��$y[l��-���S3�`�%�wU�Ԯɂ�a{�!X��oap�9��t�T�]���`מd�$2��v�0���聕��b~�`��c�P�k	C�̤.+p���}*D(�`ؚ��R(z��0��h���O�����gE��*�s�_�z�Q�I�k��9bh�း�������y+*s��̭Y�wyP��S�N�J�����r�޵�4�,�3�qo�����Y��d�C���Z{۰�S|��+��ilT�4�)�o��m�>�sa
���{����d����M꤬��N��{��\7�g� }ot?Z;��X�53!wC��4G\�<߭��,��~KԴ��v��<Q�Ê��au��J�斈*�^�v�J�\	F�0�f`d�8��=e�a:{��E!v>����p��)�G��ѡ�'��ÊF��_X�޺�¨�v�@e T�)a�p]���	�!�ޘ�$�N���(ퟦ��J��wW�a=s�pQ..�_��hE�m$M
l��w���m��e�(Vo��S:�"��A�}KR��~��vq��t9.�31n�Dg&��X�p=Qà�����9r�щF�d3�IJ�k�Y�A�����'�G�!"��$�UX+��_����0-���:9�!ÙuQ.(�̺O��Q������t�UϪ�r�հ�a�7���/��d�4�>i��Ɛƭ�|ñ#��r�-��|<��ܦ�?_�>��]\�V�U�֎�+o�7��Џl&돨����V��|��R 4R�7���
��mA_P	�k���'��ǒ�N(1B'��.S!ɜ��؛����v��.��{�@�של�o�ݬJ�����'���%-�<k>DvAz��ZW������Emdј�����_7s�}�`.��O`��D��=g���0^����enZ�1T��RO|�R�������O�-����w��Z�^^���h $��P�`�0�#�`u�F~��>�)XIq���ѳ�W�\�Ez=9���}�Y�D��p��x����P����
�4b�z�Ί��><,�k%�xW(ˏ�+#n��= ��y�
{�N�|�}m�vBx0�j��3/��:���hxt�X�~;�	�&3�>s�_��7wh*(|��5��r\;c��;XS���YU���۠���Ki�HA��Ֆ�A�h�d,�
�Ǚⷂ����voW��""Bn�xbg=p\Z��
�[JJ
!��G|�aK���}�Uu�qy4]Hz_��x�TC!Y[oD�j.j�l���qz�Opy>^3�>P�b	X:�p����cll�JO��U\(ߋLKx��<մ���S4rn4555tfePB�*/��z���I(я��_�k,X��[?&ϗ�q��&a̫�ZM��w��P7��d�Օq�Ё��Ns�����;+�'��s�kk�OWjgϲ�������^Ū��9��T_�^k����jB�����p�<���[��܌a��ϟo_S5M-,�xx^��gZ	�g�+��\?Zݔ�=�!��{�/�oG�i��~B0&bc+J@�uu?�spL՟�w�׻�����C��~o��@���:��������u�j���Cs����#ŔC�AT~gg'��[+���y(��ƾKNM%�ۼ�HZZ:�ס���3:>[��ׯ6I�	II�;N�,gO�o^O���ޜV�Y�A8W.�VY�+�ܛj���R(������deŁ���p]��dU��]�G�$�F`�t��p�Bs�����k�7��J���\t��q��q�j�C�(k�E��m��3Z^���ˋ��R��!e�%�!hi�n-�y��Ã^x�f�U�p�И�ZB��QE���5�p ��bs��b������w�!x���z�� �db�0|���,���u��D�E�4ld'hi+���k������������mfq���:,�o�^��3��
<"s�yX����/1 ��ǐ�[��y5�P��*��bM��!�XF���9�����
*��Z8��Fip6�6�5��tMm���h��!͵e �G��|��e�!�]�)!�{�E�з�8Yi#fo_�l-�.���~6��G���z#� b�ye�DDN��_�{���_��>�8�zK�,�_��FH�����ɇ\���gV�|EG��<�1���Q	)��H�������v�ɿL�T����e���
���OG�TF*>?�g����=�u�^�+g�{��#����Ys^iRÈ��B����K�Ķ4��BeO}�4�a���y���n,��S����_!Q��
J����B���K:M�f�����]}V� �����.���kk�qg�͵�O;���D����
�4�]A@ HP�Hҫ� RC��(�{G�A��A�� -t��J w�����s����ݜ���}�=�<3����Бk��Ln�Zp=�.旐�/9�oڟ���ƶV����"���2�=��$ߧrNq�9���2w�|w��ר����T��&Ӷ��MR�G7g�{,���gl��W1�X���_%z�"�����-9�`����_^ِkf��;/�s���9B�^i2�,��&�m.��hN
y��2��ry��/��ƫb�L�����o�V.��ug5�"��x�y�m��N��'�)�)���-������az�H��}��Q�Ļr���3Z��̱�g0{��	��*�V�/�u*v�����1�|{�l1��.j�ɠ�.�[�1E��æ���(���$-����=ط����k,4i�||`��3Qi��s����師��B�S�Er&Q��d}rN��	���f@�g���@)[=�?�2�ݿ�&*���+�}��Y\\,"*��j-q��n�%&Ջt`-^��o��W ���7V��ƪ������۾�HZLѰ����B����QO����Se2��><�����h����&���������S��ތ5��Q��P���-�LHi�Q�]ޗ�WA&�3Q��Hr�U([+��<մeҷ����$;�k���X�ys�a�� �b�c�.-�Lh~tݟ�t��)y����]ccc7��c��5������F�P[����~T,k�:�mu�t������[y�|�O�l���]�*�/�b�$�(��Oi�`���q��'^�e��D�-��$�q���Qjt;����`�	�G�؇���s��8H�3aTI?q����`�39�����RBɝ�L�������x��l)���*k�V���ې�O�W��L�e��8�s�K�ɫ���@�S���-(���ȃ�h���O�e$ě%?u�1a��Sv�m�cwĚ��La��X�ZkV���s�p��T��93�::����w���'�m�ȴ�4�������kWW�t���t��'~k#��=��l�cv5���ו��MT���"Sp
QśUo���a��'1�O�=����{Qk���
����7��Y�zEE�~�7a��B�aޑ![gG̈́~Y\���pe,�d��w=F�+m9�l�Oj�3����4X�mxL9�	c�������r�^
��_
���.'�Z��8��������C]{�1�<���7�D������)�Ϋw4����d�,�f�/���씙���H�Iv:.����˟��Lyeanp�⹫���y��+���1�	��je�\}�bO]����g+��Q�Q������5u��b��d��=ςPp+|=v�;S�C9U}��TX�5ex�*kc�~S6Y������W}=��ӭ.eZ���&y�sx�0r���L:�/�(H��U�^+�-�t�h�Vii�?4��(K��>c��(W�����8�ZA:eE����-*.E���3�[�M�z�uk6��d=5��]w��xP{������|�P(�w�t��5twT@�����M9��n���&cuF���ju�Y��0�k�rnM���S>!-��;DF�.˺n��ڻ{�;�5�#����{�u'���S�j�����t"A)L�;��G@�t` ���hű��o���b)��Z��jas�����R�<���5Nt]M�c�y?N���d��2��a+��Ɉ�)�|+��)���ͩ��.���\��lD�Z�[�����'Jy�o�Ve�[[�U}Bm.ȮU��g�^�3�)�f�׈��,����������!�x��ֵ�Ͼ���1��l���P��lױ;>�٩@O�˯'/'.�S7s;%U��1�P��^��c�vD�񭣘��C�˃M�������]�k�,u�o
;aC.J��~<���zÕ���������h� .���(��,ش(zU;`�3J�ZI�U���e�ƴ���{�Q�ՐLk|+A{�C���k��h$=��p������@5��{�p�U�1Z^_�'����KH�k�^teY\�u��P���i�+��g�h�^G���UCT�J��/�k��y)��6�E�'<R�za	��������]T�|Rq�����1o�֑Z��Z��-���%e[)p��#"(����JJ�`�7�u����8F��hx�}{�Z��)9^�"}h�6>�$!+mo�Y8g��l9'&6��\�o,�H��6f�,<ג2S��=�7��!(��������b�T4t�p���޿�O�+y��gf�SU�2U)-�!�NҾF-%�{��2���w����U ��*��H���Zt�|o__�f�'�`ȳݰ�^�������ԴTۣR�m5#7���z�0c��E�8׳�5�ظB~���z\�b!�c�֙a�l�ܖu-6duoxh��d������}G�=7�5E���qs�=ѽ����$7���K������)��/1�,3{e���+�,IIIrb#�m�'%�������i���ui�[;/�Bo����`���ǿ�"�&��f�}��
V��]Z�^8��9|.�sĘ�ƾ�q������m��r��˨��g3���O�v�gEEE��KŚɥ��7=>�W��-J�Fvp<���4q��m�e�\�<:�����A����M>>��s?r���g�E������k��u���Wűz��L�����(��:vj�j��f}@ژ�ԝ�^�E��	:�כ�%&}��!�UUؒ-�ћz���������	�E�O���y�2�F�W�����~ȶؤK]437	����܉�8ڙa�a��p&RD������s«��r�e��1�e������	���Q�<�f*�^�$�S��RRپ>>\����/�/��T�j��+!�|�"����#*-(t�ǚ'��#L#�kx��ƒzx��E�l���z�o�"t�L0��x�gD�&�X#"�jVPPд%$�(�������r��֝�bQAal���/���B�_�6��YT�� ���@��+��
%�1Xz�Cj<׎�Q��R�1� I�e˼�F#�<F�Tvo��f�ƅ_��|���2�-�[C���:E�ׁ����{e�+'��-!�Zl����u���>D�3���P���>]/ 8?�u��7zЇBB��s)�*-!v����i�^:���MuJ{Y���]�"�����x~�4�Т��R'�R~9� ���{Ff�ERR��������?�l�I~}�޼��4�B�*9[�0V�z�U�/�<'�\~���,�R
V.N�|���W�R���ba$S.�|����S�._߲�ކ�s]3��w'+�+�����<h-�4��|��.��gW'��q�7�s�?�p�|4���]��*���2Շ�_K�f��Z���z��h�s뱝ݻ#B�㹕p���l��������1Ny/0G�Z�Nf-�+I��sj,��¥Ug�d�J�l?G�.����,?�wEi)PD�I��ܹ
��mw�v|Qt�y���s7/��0��}���N��«V���弪L\�nf.������o8�Ǔ3Sw�ϫaO������W���mgvTU{���vJ��/���Q�S�Ҫ�2��-_3W[�b����w��V���hu�x�hXr?5"�8pg.��[���e y*������\1�/�4��k%�/#��⾩��}��GĹ�L"��><�]������+��e� �i@
���:���b*��ꇨ���Gbn���(�A6Y��i|�bv���u����A\כ�����*&E���+�q�o��?��r�70h�K<Zl"�GW�KQ�oQ�:C��*Vڟ�1�l{ܰK�.�?#p1ƽɜt>�~�Х��N�&�m�ƮYK�c9'�}a�x�k�A�^'�����~�������.������*Hdff6��qRڇ�y��֛�`�	::��i�Z��m]���X��j����5��0k	��h��L�S�+3�K���n^`��L�7�t���A%l@k�k��V�n��OgZmA�C���l�Z�(�����ȕ�yߕ���α����C>��|����Ze���9�Sq�(��˩���k��P�R^����n��p�@Ս5���KUؙ���>9M���[[�����+@�I_�����w����0\�s��HW������G��G���kp� �'�ؿM^�h������H ����uʝkq�{"�56��$:KMW	]����!a�Ȇ��_G9,�������b�A��X-��=]]k����t���x{ץk�G�a�M�;��G���U�HO�����fC!���C3iǅ���xxy�^���m�A��ee�4M���Ȟ�nd4�m@~eP>h&���t���{K4��>�/t(?��ܽ>H�Lܛ�{}�`�Lf��뛎�<)lt���n��I���z\ߘn&R� ��ܡQ���{�@�b �|��÷�Rls��V]�����f4���
��T	���*���*vZJ��xLCN+|���o)�91��62� űKo�c�K8����W�����F�a�A�m�Ɇ[R�4�(휗+}2� �*��M^+��n9<˯��Vڗq�%_��y�uq݈K/F k�D�C֋����}%�xȒ���o���eGgqX��B���W����y��Oţ/�Z�g �އl��K@�&Ox������xT^ʗ+8^��������s��zc���X6�%���P�Z�	��Ǘ�\����@H?��g��\H��\��s���L������_by�����g��t-1R(Y����R�4�m�y;��8���㸼�V�����r=�v��TO)=���6�X��\��*x8���n�cd{�۸�O����9S�4��@!7H�MG����i>{�\vM���]���u�ܶ9�5E��jk{{��JN���Ae��)�fq�Z�x��[B	le���۸�IN=�+V��x!�CA�*ЦJ�w�{�6�s�w7�-��ͬ|�%	�VLMq��4�(j��U�1�95;�ۈtť��+C��E�'���/7���Y�y%�Z3n�c���:��
9���ٳ�T�j�q�h����}���r�ͣ�!1��d�����Z���8�?���%�4All[���
�=6�����W�8�}<��4��Y�φ��s�;2�یL򳒲��P���ɺi�_�.�3&~�g���>���4a�	��_΍�\����<�'%%e6ό07��ݽ1]8Z�O�T�`V��ds��Ƿ/�)����/(Z#�e�	�x1�����c�N��r�Of� vP&�&Y���r-�_y�Ʊ؄	*X5Fڰ���|D�$O?�΄0��b+%%�����R]Ĵ]�3�h�ƈU��I0#��{ǘ+������݄���o�Ĕ��l��M"i����ʼ�X����n��:H!(��|׸�B�a�Uj����&����N����[����AK4�\�f�_�#����S����;|��w)���+5�;2�<)��Zj�>����\8�F���������KVψ�
�N�*!]f��g�V8L��Vm�z�&�$N��Qg�-�A	)9���dN�Q�-�>	��S��g^�/[�r�sȋ���8��l7)�!�^|��� [��$�y.�CU�~��}�V|�Q@��!��xГ*�|g�ۂy�ש�~6daA�H(;ؕ3��W�Yf��+7;y.,�Ը82�S�>�z#_0ao���'�N�V�?PXd�&�S�;x9��i����m����m�HI��}�Q�_JI9@�+[��/bS鱕���O�KY�|0|n���W:�]ٵ&<L�����[#E-��3��ɋ��J�s�"�Bl�GӍ�_�����>�)�=��� �Ƙ����r�k�#Oó�KVX�B��.����>��I	�����X NQ����b
����
���ι�g��'��pn�.E��,���u�����-�ԍ6�]ʲ͆��/���Tn7ݑ�w�t�L����r_&������Sz4SR�ϟ��;:~����B����GS��S�z��?��oI4�m-�QLwA P�������*>��`Q���~ 
v��0�E��0�B�J(:��}󿛬����{�,��W�ڳ���0Y���p�������>��	tC򆤸����ԃR`i)���5II���AOP���������D������E 9�c �	���99�:�A
�f/����l�y�tt7U�=r���yz�����9ہ��X�����KJ~_�JdD�20{{���W�����o�玗��#������I)9�6� ���8���>0/89IU����� }����&��4�tU�Tl#�PK   �e�X��) oj /   images/9b962a8e-14b5-4317-8666-1954827ef6fe.pngĻg\S��=�2�
��>zSzG�w�BT���	�����N@z��	��^H'z �����|_�{�?~��疳�.k�}�1TS]��������\IQ���z"�k����Hg����\I�O��ߟo?���I�Е���������:�� ����������ks"OOOk[W��N�<�.��(	Z"���d��x�m�{������O��݇D]kg`%��1�hU�O\dq5�Zl��|�M��l?���c�0*M���Z�ZwN��a��j�ߕ��b���������ad�~���ޒL���~0,�Ƈ�/�7d�|��b)���_N�;��3H�xg���c�AA⿏eri:��>GB��},��i;�w���J����S��E��ٮ����G#�%�ܨ�1T�{���''=���']|޹U��]�b�E�џ?*�������W 
�_@�O㩤0͌����g��A)Z,��m��ąO�s��V��I�k9y&�+����u���58����|������U�J�t�ر�����M��/���;T�1yD2���k�K�%�$Uf�U3�W$��B����K��"T?ϗTa�:�
m�p<k$��W�����YeZ��<[
�7.�����5.����/���y�_���L�܃A����d+�̿��!s��!s
�W�B.�@�r;Ku�&bt�����4��E�Y)!S�!��,�c�����aAX�J����e��[5y���F�,����f�i��x�d!H��y7��<�_�Mv�N�Q椽�Ѹ^y��-9f�q�~�q$�W�
^5?�]�?C��5(��`I�VZ��4[7��|���H��[��S�M�_�ߞ�x"+P�
*w�M�n,5�p�?��}���y{�|y��omj��M�z���4ŉu[_��'u��}�f��!f=�J/��do���{�+��鄩A��bKw��|�1e�&V�~��I<G��t�1[ˉ)$���]w�ޝ�.Γ�Y�"pi�s���O��S���ſ�2�Ϳ6��]�F����n4JF�y0lM�C��!�ު�(�AX�o�֮�Ue3#y����ٓ��2<�`�;�C2�Q��J ����N��c�u^��a�&I�^7 BN��pJ�G��i���q��	�j�tǉ�z*�?v�_� 5�[���W/���)��6mwƌ��%-[���8�.��'7r���xћ!'6^�h �����g��NS��%gvu�sώ��.��7'$���J�L��}�S�/�}ٞf��|�kb�W�)��ء杜�>v�zQ{P�uoQ=�����d�ꃀ��b����uM���պ�X*���`g���s���㍋�G�G]��H +K��,�	��RC�T(��3;��Wτf1j��D�!�%4[l�w&�e+�:��zI�^5x�2y�A�9���7N��e����-i�w���[���P�Ն'lE��)$�ɏ���S��0�a�!m�� �`D1�װ(\o�xoz力�׋��D�߁ԫ]tg�g؜!��C���t6j٤��� ���Z�=_���c#�_Q3��}C ��$����mD�$~�-��I����8 ��Y��3( �s���6q�\�1m�Rc�B���Wu4~��Ū��h��2��z�(|+�q���9�h޷�+9[]�TS�vW��e�Jr@rB�g���/[a�W�1Z��������DeL���O�OyD��u�ԁ%2�(�����{�F��lk��L6M]��8�z��T�B3�x����Ⴑ���gs׉ߙ-�^�6/�r�O�CV�3Z)�]s�P�!:�۟����C��9j��Pa�2��l��j�b���Ml�	��'9E�v7>�o��V�1���u*!�h��ίޕ��	2_G����v����X����D^��l�I�YH����z�����Yr�I����g�}Ӫ�a ��c�Nb�wO�ݝ?j<������Ĵ�ZN�]`�
(��3�i%_�F�s�� H�U\�fz��kw6��w���fË��9}��X�Rx��e�y�d'-�� ��!��;��JL}+�����S�{9<���a�0%��i��U%/�X%��T#��'���䡚��3V�[��)\f�3�H�y�Y<�c��j%��o���vR��F�4�=��K����,�ұ��؃��`�Dim�i��b��nNT�d|@yLV&T�-<��|�K�1��#�����;�W�s�^���]p�髀K�ـO��.���?��� C����kLLH�#N�g��oE��NF���|�e�����!����	�W1E�!G�%�^=;Z�f-2f
�36��.{6N�}�S�;��V�#�A��އ�E7Hx�"t�t�m?<_՟�?��D2AkMb����P�Odv�.r���c�"�x/��|m��A���f�8qr*�����b�u�����W3%^L��[8�Y!Z³kG�7k~ز
�:�S�)
�����l�c\A}�����L�׵�o�Ε��`,���|/��K�G]צ��h�����g���s�f,��4��e2r��Z~�>�Do��6�C|v�g�u뛳��tb�CeOw��]�c���/i�t�L�N��{�7+?�pя�Y�o �W�g���u����&
F�fLd��o^����>�_>�����Ċ�/��Y9dg41���w���:J�B�s��XG��+`�<�vp� �Ê��2�&����!,��nw�P���ك�-�|���n3�{�����w��|:�n�Ȟ��i�~ʑ���;�l�}6)R۹=z��EH4�_��W��'�5���.��A컬�l��_�p�}�����'����ض�Lz�VΥ�/����ƌ���+��J`�hZN¥'ŐS�f�M�ӱMz]Ig�Y�8f��]9M�Ư`�SR�`l���pA����\����u���M��#g�!H���Sy��fm������CO�-�����y��U�&��+@e�Ǐ"R�1�4��T{{����LZ��Z�ж/��}���#U���m����:՞��g��ɫT��k&N�詝O�#z��"{!�زw2�n�r��<8�c�]jǼU6�r��r�>�J@n�W*�U,��|�i	a����˼��oB��~|I�X6�h*k:���݆�Q�G�M��P4d�3s[p�Uk���qc���X��ں���cCs�J�x�-R��tojg:wt��f|�9=�c�a��s��J~�RWs���E{"U�G�����t��tj�*��
��1ũ)��1M���ԫ.=��T�㙫�
����q���H�-u�H�0=¹@ؿW�Y1��JK�:�"��J�\=LJ*',=�g�G_{���I�~l�b��w��G�\��Vk��=�juڡq~�˪��:w�q.��&*XUz�"�Ķ����ι~}kI
�w�2�^��>5u��?5}��%N�*�@R��}1x ���4C+�c�����i�Խ��*/��3����O/܆�7�[_��W�).~b���������72�}_0������-Zluq(���*�Cb(!���G��.8[�~��ɑ'�y�#�N)Sh0��wЦ>��� 9�` 4%�	�m8+������� ��W(��Mlg��f�z��D*�-�ӗ������>t�5t�IO�]�v_w��DA74K��u���^m�1��q�6��xp�'q=%����AP^ݘ�ݸ�nt�t���t7e�Y����^r�]n�b�f��[�¡9�o
����8^հć#n�w4��*�}n(���r���Q��U���i�����8}k㟜o�ש�>y��,�;Ѧ��b�y��]z)�����Zo��n[g4�zٚ��ܖ��i.��[8��L��1�r
&p��{��2���/���k��G�I��%0R�ۘ]� f
�}jY����9�a%�2��]�0�Q�������k|�L��&�Txlʹ>��t�&[Y�ar�}˰�����F��q���L&������;���/WdГ��Z&��N��|�d(j��-b�r�^Cֳ����ܖq��V���|҉u�:>Hf*��e��벤�YZ�3BS�����|JQ��!�6;^G�#�g	>�v����L��yºL_�,N&"�����u�Q����V@�w! �������m�*1�S*,N1�g36�B��J�=2�o����/�
��L��}H�����\��+���������"NwC���-@*�+a���&�({� �����x\!���ԖJfc�ݧ"lL�J�R4ob�.��}���I�d���d{�DB\�l[A.�k�@����0� u�D�	��y�	��	w��[��^'�r���	�ƎިC���Y��B������/���P|��t��y�d��Y���)^6�{�:v@��t$��|�-�&.r��>� �L�zGjv}�	���OgFq��?6jF���)�
��::ߝ�^*���Fz��nOn^�8��W.ǭԂ��0L�:Q�7�<�~���7���t���эh�I��?�@E�?�o���v(:�����5���󼳈UW��P��Ʃ�8��~��h��YN�r�Mi��BNW\D�m}�θ��a�c���������}�)z�l�j���-��1S�;ǣ���л-�`"���$�.�x)xi׵!�rf�:ޗ�vhVLdc2# ������qiݵn��C����7"s�#�Y������lR�+�0)�Cݷj�yK��I���TgҮ�䮇'�a�׭=Z��ўL;⸕*�����@�ƛ�~���-�-&JL�ĺ1�bC�D�r�0�%��~�g\�3���=0�o���=}JEE�ǃ�3����'�/�p""mO�6K��((;;���ar�瓼�B�r���^k�����7���?�\&FIg	|�958*��Jζ̩�GV��!��8�v7�i�P��jɯ��z��p��7}/E�A�W�y����ѭ��D8e�S���1�]t�|v��w�v.`/�Un��;�U�P����2�d�����;tH\R�4l-=l��dZ��(��{��^�-��2��(���0��0��CF���������J�--���޷�_h�M��I�ޭ���y\ ��p�*a�;z�K�G���?S�B@&r��RC˟���v�Z�$�\v^��I�܈n�;[��W'n�~�@7�> �b��4�Kdq��[�2|t����蹃^��6�JRp��@XES#���?G��:�{�*/le�W����yI�u�	�~���VXכ��
����~Үk���['���1_3kO(h��4�Wۍ�$�ac�|�>e�  Ks�����'�c�6w$_p�1���c(�����~Y�u~��i)lG��k��&w��',���B#�ё������m�u��D�!)�]� �>�Z�2�>�fM��-���d+���v�����+��(��S6�X�B����"zLycC�рLm����7�U��0_��l���~hH3��N��JD��1aP���}[z�W�^x�Rt�;��<g��2kS�V�g���W�yꞶ4v�;�\'��w?e�۱�]C��{S���17�Q�L�����	�Ļ�y��\I�y7F�)�uk����X�D7׀K��
�yQ
��ρ��rXpm[[����$|<{�ߟ��:�S- ������� Pe�'|�uF�*:�"�6��h��6��w����:��=1m�ß����-��"7AՕ���Q��/��s���ve+�/JԣM`|��f'��@����� -��͎̀����!�w���'�$�>@:= ����F�Syy�3��D�\	���C�ʒ3�� ?_�U#���g]�L�2��n�~+}��ח8_�o��a*�X5nSD�w��s���g�"��~�i��ްO�mLs���l��}�WyV=�^���(�*��c�Yy� g��'l�Cl�M��X>�U�.�\C��+B���hi	��v����{:&&�[ȭ8UsC�@�L)�P�6VV�<��Bm��y��JߑXXі�`x^Ͳ�Ӑ�~���x5Ke�޳;�F�	"��k�BGJ�,�\� ]���b.�aC�ً.��s�0��r{_��8[� P\ķ���������ʠ��+���f��k�a�ݦ��!Q�⏐
�pAMދr��k�&��%3J�7~�%��f�n���ښ��.HI�U�@`3�[���޷~���9Z������{=��۾�i�9�s����k=<�7���8����;�!�~����\g �D�筕����~^ѧ��{��"�H)l��h��O4~|�n��?��d��a��HU]�A���L�k[�]���_g5&�V�q_�|��S>g뭿��a����U�����9
���vp={��O7���u�ѯrarّ��ѓ��2[%Zmk��_O�l6-2YTD�f�W����g�+�q�w5�~8���8�nD]�V�Gv�3"9�,�M1ar}��m��E����"�{Y���Q����6�U��U�,ܒ�#���t\�dU7�`f��ҫŴ����0Om�e�:77��OC����$W��=����x��{ �X[~�2�f%�8xO�X�[��-ADV9o��D��%#�G�\�3�LR\V�c�N��}������Ís�RuY�\;2Tb�ǚ)��3��V���I��
Q��'���5���F�&
��$'8�f���A��ɄD�ۑs�I'��𻛺ƵVJ�M�?��U��Ǜ'�1Hp�<�Rݠ�U=b_d���)�Rf_�L%|�`�=�]���,�+��G��&��F;5�,�Z�I_X+q�Ln��ޙ�~�|����vT�5�S���v:�P@皂�V�>ݞI,Iٔ�"��%塡ɬXNgh5�w:]ۢ��A��*�*����Z@����H�L�;Jt� ;[ ��4m���N��6y�U���kq���7��������8��3�m?l��'ޞ���j4���g���b��s�U���97�|���`�{���2�1��]L���)�6��k,��Ї�:å�ۂ�<U\*�55F@�3Y�_\T�g DD�a���ɋ�����\^N�.	���^0�^�R�����L�c��9��S��I��}R��ӭ����iX+���~�n��˵�
�/c5pgS�r���9���e2��!�=�#��W��j������r�]|��>Y7�\V����ɪ����[��m�J����u� �r��@�1�6�1�ĦX�<��`�e,2!~d���ex�b��`�ܨu.�{�h	�2�9NN?�'�S^B���wGa���3�9��ɺ��PBo�9�ae�Z�^8�(�``��e� m央�Q�G�T�a��� ܌���Gg]0���^!���k�+�U>�kvWx���l)��&�X>��j��7��e&�<aw L������>��!���S��B�m��G��>!]��ʟ�j�o/�PQxQC
e�/`jS	?;l,07P�5��a�ѽ4���o��#P��bwȂ?[�l�q7P��'H��G@���_nشS�FR�ZJ�[v�vO��q:@��u4��8�3�4�z�f�����\[S��\YCW���0T4z�-�U��J.G�m`
m<����e~LoN4 1�����5��j�pj��#j��x9w�C#SA�����
K-�xN�.�K�i4�o��(��D��٣���K �dP��Ј��{6��@���lʞË�7K��*����@������'������:�*�mp��^���L���Td���
�u� �n{�f�j��)�;�d�4��Ƚ��6MQ4�
AO �|��\ݸ����lD��ig���o���Tk�&�S�q�ǌa_�p��Õ�\����d��aR$�buچ��]q	,ݏ��4�6�5އ555��&`�@��8>�.� ��>�N鮸i���Y2�iP����c��<���p�l��;��&Ӗ��=�	�EB�C+no��Y�ۓ�<����J���*�l��_P�P$j2&Vr62C�ѱ�m�Ĵ�d�ׯmn�~��Ͼd�Y��I�w���H����ۃ�z	ey
�xYH�5AIM�<\�J�Bi�9����SO2���J���u(���U�fC����4�]V�o��������J\xL��j���o��wg���G���tL%A�X
 ��f�-�]E%wa��lq��9�ҿ[���c�]�� 8���I(5��b}c�4����/;8덧�G�џj �~+�6��?�ߜ�,]8�Ձ������U�MTd��;F �$v/?��&t�z\�2@`q�|�?�g�.����Ϸ�Y���j&�%����yԣ�j����F�Zw��C�������c�-[
+�B�aUE�S�<~j!m¦�Wb���j�уy�K�vΎQB�_2���H�`�|mh�:�^���zA�Զ���f��Q4������|���<Wj�o#���zNm&��	ͭۻ�k�����o�x�=��N�pz:9�9Jh5�=����&H��z\�����X��1��������s�S�rkF�	K4?��c����]ߜ��˝��v\���ޙ7s�\���#
I��SSu/�7V37�f��ǣ	���	�U,|'Y��8kd?W����������+ ��6"�]o:<�]�6E���+류�I�q@h���Y���{(U-�ʤ�ؗ�.��R�C��q�s�e���"�xr��/�<X��.VΞ�6�����|����%�\
Ҿ	� ��O�����Te�X��9��%��x��녔n�i[�)���El��4�����[��u��ae
�SVSX9��<�Ǉ��,��	{n48$��K�T�G.�D{{�k�����k�mG;��F��|��2i�m��r!��N��2����.��?-�a�C�s�,�d9��y���G�r��6ڼ�>:w�:�	`��H�Y����l��#��zxdZn�Ď�y��X�:/��&���%��0��<X����RW����s�yK���L[Q��/�ϛ4�6�-_�4W��蓡B�>�ΰ��۬��O�QI7v��fKh$�be�����ٺp��z�����WA�)�����vH�h'������2�bz8�F�Y\
���wv�j+ʗ��LM��K�<d��l	�j��ى��C���&�W52�"�J"B�'�*-(��tR�����р�L���5�"�~�'UjZ��j1|9o��dT�T� F���P��`���.��e^O��Lk���w^;�>�*�=�b�����+Qn�N����Z����&#_��oV/��۩���νKZWrB�A ���w�b��I8{=I2�Bh�MM+��vu���8A�ˉ{�δƓ��!I��풴| e��U�{��Z�£+��@��o��B< ���H���K�s+��R/pn�@�-��cִ��\W:�W�x����=��e�1�g��Y1~���e�$'=~����L|�d�|�~�/����/��̘V[�kmCKe���r}s��_ӥi���+�م�Z2H����v�ϒf���g���b�V��0���H���ݠ�H`R�`9���ۏM�o�z���,U��%G\Jt[�:�Ӧѣ�e5�0�{�Oj����7OJw�u��8}D�X��(?�d&���{���`.ğ>�;��Q}�f3ͣ���&.)��#����+5.�J�A=�o��o&��,V���Uߘ��5*5i�`%��v��z�;Y���C�Nf�D��{�SV9w.u�������ĝ�����f>B���^��c�����!�n���O�*��%8�UO�������S�'��6H�,uO��rG��.]�t*����a�_8����ky��j�琎�
��7�\���/����_*� �o\ҥϊ�s���xr���!U���0��������,�`�.(���A8��H��B��*<����]2v���f�R���t����*�
wqO�F\H_��I��R�;W&�g�	Cq�,|���U&�f�=�"�݁��W13(�����=����!*�z�h�I����Cac�Ϋ�m�C��3	�Y{��@]���u���������LWZ���p��Yc��;��|@l����*�/�*VC�v��[��)Z�`�ӝ]��y���׏�ofl��e5��d)����PJ2���󰜙0���Y�Mݳ0��YQ���㟀�^b���|j888X�ZJ��&s���x�P��b!f&w��a�`��	v���}��](�q��<Sx��t�-��
��*�QU˲�]��ˊ����W@��dq�]ۇ�������N��T��ap����4a{$#��ʵ��#�XP�<$���#\@�8�-o=eT
���Ĳ�C��FNx+�+֓}�)&�M��/���8�ш+�X�����!$j�=��{�G^�_ NN�~{5���R| Zvg��	��Q�3�h.X=Lf���ߌ����lQ�=��O��ٚ�/o=���ӳY��,	�g���s���3�M;S3�*�9bS�i�>�OH����3S�Q��R%�vdw�1PX�.����oD�D���a�,�g��l��U��IF����5 ��}N�!�R�V��Չ%��c�$Se���Xy��i�}B颋m.��� d�2U�m���#�)s%�}���ˏ�O=�u~�z����=�81�$�1F�P̳267�3Se��1�,����0��'����䖅����D|�(�l�?�f6�1�����>(p�.����1E$G�<A���p$���t�����w���QNr�nAY��s�I�Q�)A���������F��i��q�H�\+�wi%9n�'qU��%_:�d鍋;W�c�?�q�5Y����k���c	۷����t5ޜ�s ����H��bH���Ÿ�.���Ƈ2�x=��zV$!�{C�r�y�� \��<��{c�_dT���	°�ժ;�py��顺��.)��םO��b̊�V�Yn�Z��0Wre#b$N�k6-�+3��?��%�*��d�!8UH]�w���z�ґ�Q�L�a��$�T�A}����E�\ �Xx����?C؁����bM@:�}����͚<�/����`d,W��(��^:�s�	i�V7�1e�\�c�l��G�
�˰𓾰&��{Ҁ�q����^�48}:���j�=���X���3�ڴ޳����:l[���w�o-]�����i�-T7f�{�t��~�M@g�L���ä������+���(�u�fվ��2[^օ���{d�Y"�0����I����!(��P���|�IҠ	���R���o�~�Q��,�4~a�c5
R$�;�{������Mռ�u�����Z5G�xE�������a�/�?W�UIy�#����@]Vb�����B�OK� �/�����6�ɺ��<x�d�@ �Q��k
�Nv.��6�Ȇ�r��t�۽؆��u�*6�YU�_fk��������C����Q+����6�ɾH��6=��Ǿ���'3rvWk��x��O�.���{,��{�G%��C{.���VF����{� :��_ʨ�J�#oPo0���[��HY\��i|(d��+��8��D'�PKk�Gٍ�jl0����2�ڱ���a�C��Z�km���&�}Z�?��v2�>���߼
~��5��g�;�#P��M	+�1���9��z$?"����΃�M��/��4�{�*.�Ѐ�����>�S���W��I�wy�r���y�^�M�K2 �NP�q��!�Th��͟X);��ʗ�H�`�<ᐾ�[�i��'f^�#�R}z�(���/kE��)7��$��ׅ<��[)�
�֍CJ֖��'��5�3�j�lPs��K��V��aO���l��YO�|��O|r�5Ua; �H�-z�a&�W�sH1�	+�#&~A)�m+�vD�%�U}��z�mN�u)�z}�l��
K=o��_�_�?�OX|��ǋ�`��ir��$�c�]���_����k#��h'���	�eS�e���nB���4�&#1Vۍ˶��I��p��ں4GIC�kc���C��c��8'��b���`k���������F���.!��N�vM�r��v�\>�Ą�7��M���w�Y�f��v}��Sb�'V���͒xp�!�2xUU����a�~V����gxX�.5�S�?����r�5~)��֪%�]{�+鼘�7Ӽ?�Z����G)iTOb������������(.Y��ŋ���P��dڬ�n��{-�	cݜ3��Z��3�:r��S��G��2#W��
��jk9nF�Qc9��lR�]�����[{Ψ�z�?���]4|p2��`EMbI5�B�+7u��fɝWР&'iֳ�7���bl�����<L�E\#h^=��B�����_��;���^Y�)`��6d����֕^����r-*�j�)��p����ϔfH}=uH-����2Ϲ�$&�Y�x}��\j�F�c?ơw�qP��nq��/���P�fs]��.����ݞ�q῁Qӿ�;'�&t���o��y���6���|��X�p�1C�އ�K���9mK�����P=���}_/�� �u(�8/ƼmNV���t�D��d�ed2M�k�0���O�N�)�ք� �ɫ�k���Q���M���js	�vU��7��b��4Ԟ���#
�Gt�B]��o�0OOx���M{_�3tw_��w�`�>v��/w�it���J�N?�2���	�Zi|�:FR�����7`Z`��?���*�Zn��F��~a����{8�X����=]��#zh>�����Ԋ���b�Yj�#�����g
.�RQkB?.����|���]p�g<�����֓�׬_	T������2b!C�E���x	�^�U��/���m�j22gՕE�����]�B?�B%��J�$�j�����,�`���}�4����<ӎ�Z���&O�k*TՈI�] ��Ӟֵ�/XA�=�[�`VN��f�"<���S���ه��b�w��`2��.�X�7�Rm�V͑�Qn����V��x�G�������o����z���|��I�?�(�ܙ��¯t��OΟ/h�ǻmZ�.���j���?���*�%�ʟ�4L�.#���RVE�s)77Y�s9����? �io���X��%�-���x;q�p�ˣA�ҋ��v)?
)᧻����Z6V0��\��;k�( �x* ;NvT��_?=��^3�xЋ�*
 (��(��m0��V�1���)�G�;�Տ<���t��'�m�����a]�|�hq^�N�	8%���Q��Ur�SF�=J1�p���H�0��m���o[5sg[�0������_���^�뽿�_RV��u��	?D��U\���_i���N�0�v3�o� ��~�ɼ�
AR�;�]�n��?���
S�N�\�
�vt.P���+K��?�_�xnb��,ȹ���b�;y��f�����Uǀ7��.���(����HQ����ôh#>b��u]L��a�/��fx��"��L��<��i�!N�e���X��2>� ��V:��3v��QB<���������A��z����!!o�X�\��_hPIE��Ѐ0��}��Gf^}��%��~�W}D�v��t����#vy�Rh�?_e�*�Uv�8Πƞⵝ&1S�6��D���n�$��F2�׳�Gقz:q9��k�3�:�}9Φ��>fmL�M@�V8̏_*U���?�;�nK^��y�-֤�-�:	h>,�w�K�Z ���}iwǡ4Q
u�K���%�"j&��t��O
�6�����v=�8���]\S�HŔ��[xzڂ��[ג�H�$?�Hz+��$����÷�}yt���WC����ؾf�^E�+��Ÿ�j��d���i�]�I/j:>�H�����3�B�a?���ۇ/z�k�:M����N}'���6�<�M{�H���x���.;B/�r"��l������O�c�/�H5OqzJ;�|�bSN��#��0ʺ����z}3�6Y��y���\��:�L�Ld�O__j\W����"WWwwrt�"��3�B�����_V���bV�Rb�Ѽ����)����az,[]`���s�}��$>~E�R�=��=3�޴���/~V��e�g�F>��]��'�MM���Y�|����^ѧ�Yeoʸ:iA}l�OO���~�uB�9_�ڊ
�r����I����ݐ�<��'�w�n��?���=�}�U���EH�%^�D�4-L��NS�%�Dg�T~��6���b��rl�ê1]����R�5/G�#�O���B��vy/��K���ϓ�|+���S65m�!�37�S���S�,�3z�
4p�Q�]��!�o���1��-n�IW)�g��'�|���'������{<��W�U'���K�1���k���kc By���� ���KW��ge[ճW����=�WQ�e�M����Ǽ'�Q��S�����mUe���@�+��ѭл俆�㲲�߸qC�g�q�h��o�ݏ�%��Q}.�T{�
�6�R��|�yk#1#����c�W����.f���Qr~�����}w;�n��\$���=�*��`�2���C�-��x�:)OjiTd�"�>,�}�_H�����p��|�������~V8o�6�^�u��ߵ9�~�
m�=�Xn�Pm��q2xp��h�霺�t�-��}_�}<;"�W��$�bl�q��-�E�dcs�rb`\�󮔺����8���^B�f�.�Ul�,�>�����{���\�ԛ���U�%=Î�`w�zGH��=����8\�2�?cgz�Nã�tx���_i(��ݩ��g�S�� �τ�+�;���P�	n]�ҧ_��6N�9a)!�mu���k��{ɾQK���ڗȑ��DP���#��I�^��b���T�{�Q��[ʥΟK�d��	�h�?���5T{,L	�N�GG~�brS�\��w�xyҼ�_�����F�u��4~�	W�A>�����R)�_ZM|Y���x��D��4��C���N�>�S�ӛ���.���wo'�<[��|֥]��ǁ���<M=�[)�ܙ��.4`L|�N���U��-�Z�Bҹ:{�TGa|�e��������vά�])�:]r�p��3.3�3u=>� ��{_,0����&fͻ˞��&%�/�����!��������D��o��a���)���q���j4����	���l�u�$fZ�_�+���eRW�|�������0�����sc	��Gb&g�q��3�t�򛿼�Wi�7�E�b��$��;���r�U�b��{�*Skrپ\�m��i�u�.'>�0�b	����',>�0�E6�|W���6�P��#�[�%4�O����yX�����2>k�D�<�����uўs�
?�.��-�����t>x�h��rҴ��a�f�)HY�o���;�
ϑx"U�^Ys�H�;�-����C�<Ðk�B\VKF�Ya�]j�u��t+��H1|��i�<v$�]4��S��U�P�9WH�?sn������5�_����bO��~�n�r��jF?�_p�`ۈ0i,w���`[%�����������r�vڤ��y7F.�Ky�N?��c;�^��D����<�� �k�t��}gZ|
���vv�8����߅"���N�_�^��b4j.42��c7h��CL5��K;�ɣ8�w?�u;btK}*��O)\цBu�c��cz�o*N\�ku�������3��F4�?)���ԇM�f�D��O润��')>ʴ�x{5���뫍W�4��nL?�tq��#�6�i�xy���49�}pP��^�+f?]#u\���s��a�1R��'����x�~ay",�e��g̶�'���;[�S��{Mo�ɀ�df'���C�\ӆ}J7�����Ơ){��[߲l)4�s��'��)��UA��ύ@��JAb
����b�
2�ѓ����q�:oi^��y%���q�V���3�Xv�n�^��_��-�1�!���͸��^�P���e��V����n)(�r��w�k]|t�mdP��>/X74B[;ܾ���	@� z�z.Df�}݁Q���n��IA�Lg;�����0܀�9�w�W�X��%#jv������C�aS\�f�������hi(ɯ�Q�5��6$)4�|~��su}r����Z���<r������י-g��F��_B;v20�ߚlK��E
>.�wS��?}�,� :0Z�}4�� �\��)>�o������q�㤥U���<�fX��¨�K��[r��S꘥�ƶ+-��1:�s}����h�(>����1��P'��wa�s�����q-�JӍ��uy�t8���$HX��x�P�o�7�k�U*��t)5�o=�#���Uǘ{������^dOB`n�����3\�� �ڶ�uZ�v������9���c���w��Mn�
�J͸����]܆
��^��7��L���]�f���n���C�[��
���!K�����C�y�|]|�������ѩ�z�5�.�ů5]̆w�)��[�xa��&i�[=����vW��[�ǔ)�{�LX�������\��M{�_�=�sx����F����5��!��]�ݤ�>S~�K^��u3r69��5ɫ6�E=����mv�[r��V+#1_#7�����J�1�,�UFD�ȳ8�ͨgs���=&&�}|�9�w;�Ь�ƽ�A��hR�K-�n���E����,���Em��e͘O�>P����{�Ze��?���q�<���(���f�q0�KV��Q2�����]1'3��K24������$�*6�c"V��\�SέkG�-wwhQӒ�����xX4�,��V���Ӎ��Am^��D���_yVj����}��O[,��1%�@q��Ɩ�Aa��Q_�����y�;~�_,
/�(8�|@`7L��PW��@��;&w��^t#���,��<(��h(G?4y
�7����Lb�I��S�7��(�_+Z���F�0\�ch���z�xc�=���k�$���k�����&�A�CB���A������S	��;�����Y�ߢ���;���0�����\׉*�ݒ��ް⛹6gv���5D�bO�!OҜB�߯�ԐT�B�\߽�l�ȢW�[�Q8���Zk].�p� ���\"�G|Q>~��s���C���Ć.�tD��;����.t����\|������d%N2��4����WxG��]�7B�_���4~���ax���!��BZF�}U#����wϊ7ڊ��s��wM��[NԵ(ԤiT_��4�$���Cr;����b�W�������B���?m�/�{��'Pܕ6��~e�H��{�۟_��L�Gpۂ�Z[��z�YD µz�hT㲷]���b�v�Ma�T�M�9���C��C�@��c��J�KY��yH��x��-�h�\����˒��m�8�r&����~�ގ�j�G�*�d�qB��'^޺�M�X�y�f�Jg���-y�l��5��_���UxU��9M<�	�f��c�4���I�V�!V����`��"�B>ka�-������%LȬ�h�S`b51ӥ�y�7;�FZ\�
�#.�S��Q2�� Y�k�>���@�E�����__���}.���Z��{+�:��
!W���͙�(�r�Z�0�^J�����/\[P��h�lR?M�
ZB䑬9��8Y�ۚ��w}��E>�3����x�8�81��wQnn�i䷱u�����z޵�3�Bp�Z\��e�RP�0�tw���8�y�t���K����7 G����x����)�p��B�q� g�;������������Rg��7�w*�]��!���?��E	_��t���j|R���	��q^�6o��SΘm�5��r�(<M`�o�s�r�!�9&6��N����+�{Ƃ��K��N��Y��5�CfL��Θ�G������b��&��]������qO6��GƧ����e���U�ϕX\��>R���p�NW$M��T������>���ړ��L��@؅�d$���Δ�Ҥ:W\Y�4��m�v�|`�[�l�is��)��*�^�����+x���%<%g��{����D	v����Y��5!���Vk|>��c�?�q�J�I�q쩕�㶉%���������^�*a5h֨}u��)k�yc����0kv������ <�$-8�~��پ�9ލ@or�8�fCH*�l�]������`���1+L�xk��M��u�o����.����?���8��w��m��*.�k��	��[*�*R�������v���bv�Lm\�v�	��熥����wϖ�ֽ�gZ-�M&x��*�̹�9m�e�.Q��$��l4�Up<v�f�4ġ�"_F���-�)v֑2�C���/,��0�������zRy�ɩh�6'\5�U�V����IV��!��@�����l����Y$+��`�ݪ���{�(M��Ϙw�wk��ri
��~��K�����\���T�����v�cf����e`��D�\�5�I��z�������8�{�co,E]�<��o����S�X��]_%�_���$����D��f���̂�L�` ��?��з�����S\�d��n���ߛ� Y����*6h@/�{m�-!J��~�
5l����g�m��ւ�c�7��[|&���ה�isC^I���f���}�#�hHVr�1w��zgf�(Y����5uUf����K���q�K����u7n"�V��}y�y�}!�'��������4��p-wخq7ܬ�S��&އ]�UP�~
I���x�jC3�z'��y"9&�Lb��e�V]�]�

���$(l]Pm�ē*t����sw�ur���(+W���M��*|.KMQL�@H�ztw7R��j���mӹ��Uƹ+�K�|t
@��t ;��,'� �n��2ŬKZ�kL�=��th�L��\嶕tt������%[�������VnR,�'�q�)�̟���u(���b�/�����sr�U_K�(��~3*1�z�v��l��c�s����o�|6)�~a<�Z�F¤������0����Q��3����鷙ߪ�1�(���A~��B>�"�~2�[.onU���;~\ƭ���u�Ga��l)d8��ψ�I�Pۖt���\�3;����r���vb8m�7*����Bzi�>�4�Ĺ	�65����hZ�AZ�ڑ�#����ר��n�KJQ���/ú�1O�'F���!������ �781,��.y���F��:S�"(����8>�����''��-��3��Jv"	�k�ר�֗6�.Y�7�>/E�N�Cg�&��9)M�h����L��[e5���q����?�F! �<�g��c⡸c;>Nd|�:R��x��"�+Y
�	kƬ!�����k��n�޵����-�?�;�@�ԭ��k3�x�ѻ>��u����b"Ԩ?��q�3H:rݷ�upq��È�����x���u�`{��`���q�:���he��+�Ն�,u��c5�,��US*�Ō�=�r�0��L���љ�N�֮��/�o�"����� ^f�]�q�-f�tl���5�� CM��M�NET�Q��T|#c���@FN�|4�O7��QDDDp��gL���=��gޛ�I�ȵ"7a������%aI��2��O6���gغ����a;�U�9���Q̏If̋��|���n#�}�Fϰ�%W]��m,U\���׿�������mV@O[��é���g�����D��D�wEBӿ�/�`��A�G������K8PgS�(�}��)��..�Ws�^������[��s*��q.[�����	����ݮ�b�cB��Ҋ	�>6����]ە$���N�[�Ǽqm4�#0�S��Y�ed�44�rhY���*�"2;���	�Ф������Cea�}�aRO��a�0�F��:X?�s��R�?i^�9�����@
,{$�z������S��rDiހ(�D���50w����N%�hE2@g��2Эwa�!�n�wΟ/	eu�ܹ��_��O�+�cBvU���/��1ש�_�;�� ��<d���/����g�V���Xr���&���У�������M	�6D���.��ll0��C{�?竭b҅���G��-7:�4�?u����S�ɷ����HQ� ʄx�|Z&u$EY�TN}ϰ�CRB��]̬�ٵ|�&lw�vK�S�6�k�zʁ�r��1vG��eҘ!T��ӑ�ɞ3����Q=��!B�nZ��vZ~bL�ro�q�v]]]$����3���M^%��{X��v�������)���k���}/��z�G�Z�4fu�p���72�]��/ ��'�Xu#3�P�)/q7�6�"k*E5��/p���Gb���9�y'~IE}���:X���ڨ����;��X�W��f�p�ՙ{~rZIӷU�j��)�J51�;mo\o��R2�Y�{�xR�V�����d�YWiQ��vZ���F�]頃�UB)��ue�m���!ϚC!X9Z��3c�y�?;�r��;4���o�gN��ܔ2�T��?63���-uBu�����*��mG�����r���
��e6��)ϑٴ����ǂ�F����|���]8��%`K�%��ђ[�O�V���^'���8���w �J��Ȧ��3*��@�S������RD���� �˒6+u�����T@�%2�YC4\M��񢢖IJ��C��\��e5a��,q��]�{f������&=�����*\�/�1y������Nx�sVjZ�:2a"����A��ba���|����� � ��UQYp����r�������S���[�.2b1��;e�M��{q��z=ߟ�a�l��*��^^���׶Kx9Ԉ���W����$�������������KҶ���M+�����.��p:�&\o��e�?�����|1�?���A�|��(�ZP[��P#hځ�c_���ٌ���ռ��a+���ֲ�?��!<ɋU����D����Ђ��p˛����kt�a�ㆵʤ��R�,��H�	��Z��8����g)�)���JOx�P���n1��ف&�$)Vof6��+�A܎�?��|�P�2���ԋ+�n�Kˊ�^��/�_�j�}�S!'P!�Xϟp)�tw�Q��Cx�S�d�j$��i���㝺�h��N��� �Y������ۏ�m,�a.=��N<�XЌ0�54�}����{�L6�І�Q�^_M�\Z׿$|��;}��N�0C��,^͋�k�C zgW���5�)�j���fl-$Z3y�(tFT��k���!�h�2&{�9-2�����1'C�CE��u�|��gE��x2	"�J)���u��Ξ��;C�Y��{'|l={�,�������%7�Q�c#˽F�9cw���kɅR��/��!Rsoǹ�/�&ٳ��!\��X�#��f,z�s���/�Y���6�5u/:�[4�,�����E��-�.��d��e�J[�ߓ��܂^b��O������:y:���O�OgU�#���f���4��"�݂�|�|�7Vi���w.`6!߫�rl�m��賬�{�bI��"sB�y�hȆ$�?�����"(�޼TBA]`�X��/���,b�	=�:iq5���c��hږ I���y^� ��)�}�^���?���L^��zv0�z�DN�<{9vv��Y���u�aP�ƀ���tdѝ�1��ތ5�(\��?�h�C3g�sM�$��C?a���
��|��hG����{߿
���������w�w�fo7�<�U��d=~�r�V6�i�� �V�c�j�^#�#�C�
�ʑeJ2�r&����n���1�'`��z,]��A�a���5ݜs^U-|_�G��b�p��y)��l�4�&�B2�iQ����9}!pS���O��=�Q���Xn�D��,��o�z�[�]TRs>����z��/U�����+ދ�>�������ן�8�ޙIƸPK,�3P�#�1�m�i��=?�H���"�lXC�O��R�x��8�����v�_���<���:<I-��2J��^e�(�O:a��;$8�:�p�:h�+��<o�C:f�,���:W��;a�t]I#���A��{C�/��й\mnY"��0w[: ?�s}�9�,����.J/	����%����ӵ0\��WN״��ǿ�^q�6;D��Y���/�9����>q�R�����y�UJl9[���R�B�L��X�~%o�Pgi�t���;{Є	�O%nud�ʲdn��6iC'�c/��n��g�&^}_������8�/&���(X�����2�H�Ȼ\�O)����y�1y�|���C"��eq�L�5S�������.�����?yx�Qq���h��d�Ui6p]N�mQd��o_1z����+�vYJ�0�u�[�i����6<)���G�2v���� ��`2O�ڃ���bÎW� �F�y��&�t��DP��c��Q~2�rDkb�͞^gy�Г4Ѝ�*���'�[�"�����G�����@=���܌��D��6uT�����z�v��W�>��_�$���IY�_�~�P���>`�u�p\����&�v����%ܶÇw .�|̃9�~�cBw��U6|�,�a��ئXWx�f���(��>݄�gOl�c�wO����ݮ�&QaEY�l�!��k��?[u+O�A����Vv���%C��Y���'���1AA���^$%{�W`���sR� 6���hpm���H�m:����j�-�j��?���dz�;�#��|�j��ZAp�!�FB���z��3�
�
ae��fUb�z9�b������S�cd!ۛ`���<�v��=��g�#�.�n�f[�OΙ7u�G�f�.��#x��=��������&�*�+ⴠa�opa�,Kp�E��m��ߴr<��8r r�SY�\��tn�����7��v�@���~�_�4�����֊<���3̒��WPN��'1c4
1��TҎP�Vf�]��o�'-;�gw�p�с��|��_�nY�}0~hRme����ѴHڢ�4� �ǭ0~{H��/�|1a�X/��(��T�I�s � �
1?�k=04i@����]~ƚ�n�,y۾/t�V�f6�.<��_a������-�z2��5���SI�Zx�z���L%�0Zx��%��F<���;��9���� ĩq��J=P:K�$�|V�b��z�6v}%�ni���X '�~Bp�.��'{��e.ᡝ��{|���e��e)3�x��SY����HWb�u^*��|mJ/��ǣ빅�53T��cc"�Y�RQ�!�0��t�!�-��<b�"�]0��_.�9��^�֯'��$c�^�u$��)l?�IN�5�?��.M�S-��ȣ7��Y�H(��9�01���M��:	�c�����%��Ҙ�h������a=� �[��߽l}%f�(kF�q��P�hq��f{. �M��d��"|- �/�k���-Ccq����(h���W�A����`(Pvu-B�a�k�Hxۻx 	_��+<2B��ٿХ���"G,������>��n�k�ׄ�*�ί�0���U�0�dwz�BH�?�-j#��rr���/�C���}�&{�㵡c;hB�	��tȣ���0a���\f�L�܎�Ƈf�A:�=;=3�������>�4�9�.fgl"�f�x��賛o�ۙ�F�~��-J��F�>�6	���T�����B�4n<$�_=+YF��\GxN�L����pUPЁ����p�����>~�8|�j�,L���~�^aS4YƆ�����'�֡�Dg��3�WHX�^����Y3�[n��1�"n#+�Z��׎��H�(��d�dYfb��2	��&��u���Ls�i��1)Vzd�2�s��d��/�>͸ل���r�0��z�������������F�9�5P�~ʟ%&��{р�{�Ӣ�˥}��~�4�u�8tI�U$����~�m+�-�� òh�/�<.1)���JT���L�P��|gRAv����m���"�m:x.l�B$b4:��t��x^�K�	q��]>�Z颎�/w�g����̩U)���Ƨ#�U�17R��Loj��/mz��YG�������\/�N.����ӻ۝����K������zOd������￉�%�M}�Q�p�O/�k�����A��u�6o�g����~T�a�N�VI�b��"�Od;�Ϯ� �w�A�G��d�����/��ߠ�F2IA{��V�2�n���jtzU�{8*�2������iK�%J}���{2�{g�#�@u܋�/�'���)s���d-����.����V�д�����ZM�9!<:P��t�>=�w'����A��P�� �D����R���d�k�
��31�ܸ7�"c�/�G��TbĬ*m^�R�}y^��LL��f�'K�И�94�P��"�\��j�O�_�>��a��tbJƄ� ��Ij7�t��@�ko;�pZ٢�6�*56$�����*�U5�|�O�o���5��m\���<��s�5��n�?2�Ni����EG��h}�|�����3�)A�/Q���Ң>���6 �l�tx�1$�}������c��IsL&H�A�"Hj��5�7&��o7J;.��;q���M�2ǧ��{�USB��'�O�)� �L�Љs�ۓ7�I�����d=�.�d�����5�c����ِc��c�7�8�Kē8�\}�����s�ګdA5`���8�c?���>�cxJ�s�6��e"�_�$��ޕ����Q�Z
8u��Z�'-��J�#z{%S*�0����M���ӕ�/�6�4wuf�툦s@)I��/�{�	�)�z2�S�j�^��d��\~��A: ��$ʺ��׹��tX���l ~�]��\�}F� �ǚt��6�;�V�xED��8%��g(�Y�Puul�S�������&8�ݜm�2�0�N�vm"�V,���r�L��u��]�Ѿ�&�\�ox�O���Vj_�|k����$	'E[�$���@<�E� ��8���H6ϕBl==���O ���I+[�LAG���s�=��;��R�	p�f\���_�k4a����bu����M��6}~M<Zo��T *L����ex���gT|<+&�v���-��(��0n���$����W��"%�'1~I��bB�ܑ��/Jb�N/h�ܭ��˿�uzˊ�uS�!0qh�i&f�"N��=��5H��K��6a��B��=����u�I�͐!��X8N�p�ȳy���!ȋ�Ȅ �
)44�&?�c���z����+�7��.�y�c�x�� ��j�����H���5vu�t��0\��\�5�_p�,4U�l�P��t
���(Y�1��{��C�S�Ab�G��5{���͑�1�r���$�'Lں$�b��s�v�a���H{y��/7R3�k���ٸ���>R,a�M�8#un�D�Ӳ)ta�-, 9�:0�����U\ܧ�:��C%���M?�$M\?i����u�˛�{wD܇-���C����giX������v�Mޑ�GC�����2%�W��m�G��XnaGiޚI&�b��2^vE&�P�r�dn�A��":�u�gJ�f���q	���q��.~��fQ���ĲTZ�r��e.Ј�LB�e��Tv�C���7��ں0���|=��s���.�.$E��T��z��vӕ~�����q�=��A��v1E��[�g��\�&�̐6	F�_���Y�Bs4{/"|�x+5��R��*�!B�4�Q��l1aP�s�>@<�����^S�gS˔�TH�cD,�'�ٙ��^��ۿ�r/;�?v%	�a��Ļ��t_�z�^�E�%����+��\��'�
1�JN�R�����Ј���o���yqWG�&� �ԥL��)7[�g���P9�k���'�ع]��6R��H؀:\VD��s�` �[D+�+ށxc_:.^�jAPƅ��$��*h܁,{� Us�W�u�-�V�~�!q����G�N��{�9	h���u�ϕW*��YHrH�m�PU�I2�}���^6��m�9��T/!����o��=�0���bb7C�����j�� u��lO�3\!��M� O3uu\g����d _��O�P
��40���&���9B�P ��w����㦃���R�|{�^Ts�qb�CF�B%z�_h��1R6�O������OH��3g���1]WPx�n�JLsH����Bs��[��/~��X ]�L��<� �0^��vk����[�3��(���R��E��}^VCYi����c����N��I�(���`߬'eX�FB������m�sm��*��ݟ+�Cʃ��uSG����S��q���_�L{�����ڸ�["�ڤg�=½=��~�Ed���J�/i�ArT�_�Z34Dθ��:e��8w,ͬj�AN��p�_.�Q�㊾6q�,s9����}�>�
KOW��v C��*Ѫ�Z1"p�KK����Xz|v�����A(qݒ���T����o" ,����r�;���$$R�T��4� o��IxD�u�2�Um��ԗX+���������fP(S�)�e=�:�P�sqK��K��vO\*���#�k>�(�X X�h�?=|��O���\<��ת8����М��.�D��fV=CS����e[��e�ӡ�	���j���b��y��[�MD2V�^�����yS��-�R�V�oS�jD$���R������q�s��	�ԉ���:0.��b�\�OK�9�Z��ؖ��'�F�R���N4}�RtS�d�.tiGS����~��v�Jf��=s;��!Y/o[�����=�l���n�C7�W#V���U��Rn�l�W�+e���(1���2�ٕw9��"���V�V%1��!ʯԚ�k�A:�%j�g��J3w�@����a�5��ް1�2/�1���g�ʹ�.�KLKl�drKg1�`詸TL�D5�M��᫺��&D�&�m�g���뜀(���L�4QJ:;!���|�F��6k�d���IF閂H �'R�p��;�#ƪD�����6#7Z67��l68�y�\��F��Y[�~W��l�)<�V�9c��3}IL�w��R��� b^"pfs���Ȳ(�j~7��XѠ7OkRydP��F-����g��Z�	��<�K+_��s��av��3'6��X-���c&�ٺ�o����ς���������'��y�\�@h5��Gp.>����lO-W諴~	A.TMWπ9M��Q�yU
�%������N�+S�g�	��$s=FH@~���(+P5���8��|U���?�_*�0n�����8$�����-@��$��@S�����}�e��ˠD;ٴ턄-{�����1��M��GtK �U��%����h�
I�M�u�\d'���3Z*`C�܁T�j�%�&��܇��Yf���;�9.$oE����gR<-�}���b���W �c*(�rE�zH�r7�팍�"y�`��,���%/���I��:zv���r���?$2�6c���h�w��=
���~|'�'P�9<��]�.�O�}7�|}����̄�v"���Y�LO�J��i�����b��lL��۰�NH/�MH�GW�>�{#�G�| �;V��.��BqA��Ͳ.\��B�%9�����*f4�8�8�!3�V���p�ӧ��HHrkI�2������҂�NCۛ_w��xW6�$�3$v�ǩ��֤�bq�%!1ŽWw���Sc��� ��n�G�#veDl�縋��P��2�/ӝ*���EQ���TH *Q���C��
�XL���@QI35)�q��,���,v���C�:����Ͽ��܃��`����8p�+�tsm�f��b֦j�D�&lS��'K��MU�ޅ�rUWk�5m&��4��-9즾�oι�H�Lzh߮�E���K���CPVu�z�JG��F4�a����,q�����'�צX=�d�?�OvCY������8ֳ�6��e�~�n��A�����M���>��v���啊��SHy�Z�̈���C��!�g�KT�<%����(��I1Զ�o����˸!�4D�f�):0�(�b�*��W(C��9��f[5��J1�p�Q��Ыk���JZ��]�g2ޚF=�<���ް��4���Eڈ��'��7{��w�D�O~���x�M[��0�囩`�>�+��"�c>W�2�v�c�k��3�J��Y�� D���Q��  �ާĦ}��\��m6�`Ӽ�V^� �1�D�g�ȳȦ��+<x�(���N���W�gKR,0�d�멏���r�mP����q��.C�z�hX{3Q!R�Ik�-�<��`��Ξ�>W��5ڤ�:��˥+��U:���pħGj&;$�#^���I��^+Nr'�����Bu������o"X[x�h�iu�8̒b�eBu.�^I�k���?[h����J0�o:��h�:D;@�S �k�9�Ci5U^�D�ӻ����R�qɆ����ܽ7��\[��a��E�^<�Rj�.�u7pٌYV���mL?�z���aw�{J%Y��_��;?f�����@˧�+���uF1O����|�g!:-X���2ESr~a����.s1Ze�k�ͬuC�^�&l���+�^���Z�X]�<���D`�X^��ћbw��{�$s��9 M�xAD��~��(���)�QJ����o�
�Ǹ0����>d�E�W8�7M��#��2idq18�)�k��(��x������V: �0 4tC\�
e9R'�{I2X��"��𑠗.���"
1�a%���Lt�/P8���p�w��@N���n(ԍ��5�ڞ0�z���3	�$D�����4���Q��҃��o���w3kC�Ó����6S����jJF/�A�ɞF��=\K�Gn�G�"%�W^Gb���]<�W ���lP��F�zs��bi��e8V~��Jt��y(����p��l�t��+���Ѷ�_�k�IS&O�� �uȦ�I{��2�Nj��LS��+���W�q�\G�J��I��99�6�{�C79��&|����������/Q�9ċԂ�!Z)m�/K�xe�8Q�%��%ҺĹ�!Wx�ʴ�
8��J�=���%���h(K(��2,J�Z������\K��4���_},u/VV��!	�G�ͬ�����8] ��f�e(��P76d�Z' R[PҪ�D�X�J'�KA�\w*���+�\�@�l�\�SϻZ�/�8b;���Y���?�����,��(�R*K�6\�79�m�Glv$i!�����5�bȿ�(��GKD�{�UQ>�1Gl����<�z�"k'����i����p%NP���j���dL�RG���[�(�oXֳ�����`�6�>��V�l*m����D��J7��2�ye
X6:L	��J;=-�b��E�'����}�t�/M F����2��z�8'�Y1w5+�\����F�|G�N�"ҩB��f*�o ��P?�/�,;y@����Vڡx�V�.�]�ZY�G���^�#P�F�pL�$oI�;Mq� eɚ>6�s�跞���B?D����@\	����P��V�Bօ;&
��8|�T�?.r��o�j�m���4N�&��R��νHO� �
7��*X�lN=�
<���'�z�
�^��$w��Sˋ��D]ڼ��P��?�,Gm�;�0��-� ;��(<Ѩ�aL�J[���^��᫳*"z'�9am�.<i��l�o&x�;s@��{X-�6G,h�}w���d���Y�O�(D��fd��v-��1����!'}�P�ۂ�2W���s4�C+"PB��Y_�`i_"}Tv5I�@<���=J%��b^F`�R��dQr�Ĭ�U��^�5�r��]IW�S���v�I��{�� &��8����v�*cD��00� T(��X>@a3�v4#���KU�<��/u�����i4��"�3&��Dm���[i�g�ތ��G��3��i0
��7L�)�М���y�!��\��Z]i��b�����v׎��ܶ���C}X�:�^N�&3�@��uawyƅ�M�*��(w�]2��YTP$+��cΖ������\������]���	V@9t���eĿ���I%�RD!���>҃����?���V��>T���vT�R����0t���#��aj��X-b��8C��X�<W�}�n� A>+�Ysj��m�Uz��$ҡa�a����l��vh`з�����X�K���u�W6
&���y���M1x�.
�� (iQh8����D%i�lxi�L�n��6qy�n��^o�<�a�qA%	�
`�e~�����:�BN�K�NP4�����^�>�EӾR�ajL�s�����S4q�Bs�&�~�g��^�<�K�T���s�/�r�����aQ��0��3M�Y�^�e;��F��v[�^���Ox���q�s�l�}�4W�/�>0�p�d����2�@r���vO(4�
�|%�mdm\�;���Ck&�z��K�55�w��]�5�AP��`���7 ަ��E.�)y%Z����Q�Ʉ]oH�h%�D<3ŉU3��<O:��C�h���3�.aJw��z�s�����<٣DpLQ}���B�k٨���+W��������y�.� �q���<)�a+�y�dC�S#V�l8� �i��To9:N	l_���_�����4S� Q������1f��ex��%ۭ	��{�IXN/��1�q�"U�E�e��˚yc"�uZJ9'h��a���x3��۔�aG�L� ��ױբ�1�[Է;D���;*C��2�WUk-fM�#U��'��:H��w:�5��29���z�%�(����dSݦ��%�%z��n��� ���6�n�dufL�	�X�?gl�O��V3E?[������4/3��:<0,�l�ʞ�/�@�NP�I�-ul�L^��=dS�Z1�to"/��)����:G1��	&Yd?��bGA����8!z)
�Ue�8�%�9#��^��Qu���Q)����/~��	A!�DN�W�bk-.�[ΑX���j�&���h�E*Ќ�W��ѦG�ĵd�	���%B�D(�O�����r\�����I��%�K�RF�*�m��b��.,h�i��MJD
4�䎴V'�mp�=<b��wP�Jw����?�l1�ķ����3�?d�9kaT
	յ~P W�ɶ�ȓ d�� It������.I��3y&2"�v2�]g������M9�L��q�!=P��8bK��O.�����d�C^�o�60� ']�P��W�WI3ީҐ�mg ^��J��[�r�3ڽ��kd(��o|�$��}%F[�1��:'��^�$S:���}��@�^Y���������&�x桅��r�T��	mDI�J������nhiw��	���9ίJe�x��ퟺ��p^F6l�b��beS '�щ������?Y,�M�4���j��
00�v5�p1�����R�։�������ҥ���@�s�Tzi6�g��b��+���ήf��;��$-,�c*�޻,�]��v��%����B�h;�c��lp��ݗ t�z�R��k����Ab4Y��I	d_��^ﰱ���F�
�n���	�8������.!��g_I��\�Z���2� ���)Cwō�*\G�.)�ֻ��k���o�GF�D:Y��ը���Ȩ�BNm��Qye���)ۯ��U�P�%қ���u���-a�,�2J.�1�:��p�m�K萲�x��F\?|��L���j"����"��6Ľ7���皎��_��}[��t��M<ν$u�����ZnrHY�/=F�k"b{%QF�&\�y���Ɉt���+�a�^���"�@���כ���vX<�����<�����K;d�@�oY��<i�W((!��$���6��I"l�b�?��g��j1��\F�"��$~�#���O=K�5�ѽ%kV�iޟ��Y����z�ϫBE�jO|��$���X�S\OM6�^�Ĺ���?����r��4��_���RK�� OO3PB�d� �|m��~��#��#(IP���ܯq�FfB��'�l�cAf��)�_�9�2�Пi���6��YZ�@�g�������+�ӕwj�'�h�7\��;�3��Cv�+)f)��TBP	R���$ϭ2�t�MUV`�#�+	��)�T���/�ȹt.?,h�L�p�Z�A�L�'Dǝ�}c���+��j�*�w�DH�Z{R3�_�Tl��o���ʡ]Y_,�5E�~E,3�2���������n7W�Dw�/�0謾��"t,8B�S;��m�z�ys�M^)�5�E��M�4�/S��^<8a���pE�Z�֭.%�ac�;:�U�
���C�ZYH��Q�Rp�i^��H�1Z����֖.u���C�ˮ_Y�ב��f�+m<[���Ԇ��lk��u��K�$(��Ї�M�		�����Z��d�@2��W�TYt�W
FhxΘ�8�Ui��#����؎շZ���i�-�1D����sZ1ąm&46�g(�WkiWU��hA�N�}��x}��@���cD�����j~�].��vzL�5y�礪 ��Ǘ��H[ۀ�o�pFYG˶ėrn:^�lY&���Oj��?��!N�t�[��N����p��w�������K��]��D>�!��#jX�&���V!w�����\$�Tm���B�U�G��D�|q�k�C�j-J�%-m�W�#�k��~���H�_Q19�-�%Z9.0~�G�YQ��*8ME\��"����Q��b�C�I�q���+�Ͷkt:�ǿ���c	S��� �_���#�'�Y�B���Q<_�.IihƼZ:�i4O�E�-�-�okp��[A�/a���)~X���z�7����^�^{?����V`E2-�ۣ	�C�����,���ղв�#���+��� ����Mf�\��a�o�{�F9[Uir�4�Md�����A��*���\ӱ'FB�2�_�S�z��PF�&�O�������g8�L&��"T<���Ys��9�P$D���ANf���bk�Y��6�l�e�;�Qz+�Q;�4���@��0y��G�\V۠�JK����݉ɻ���Բr�&L{/R}K��b����T�ԕ��"�l���?2�N�>�(�������|�汉M0�D�\<���HF����*������C��'�y?�3�ѴQ�ho�㵁�n"J� ���W�����T��=�꙼��a�}�s��ى�e6���ӕ�$l����Nh&وF�fz����L%&k��6?�sgHg�	9˴��WE0�l����t��/=��A��i��n��y�dB��1i�(�9�����Fq�Z����zӾ���!W���w݆D�3nA�,�
�R�n��^��\k��t�1n2(�r-�����Roqy�R�gO�mk�!�N�Qn��n�ٳe�_�<�
5�T�������=P�'^��(k_�m�l�ƐU�� �
S��i\Yt���K�&�L�:v�/�B�4k��}��a������L��B�R׺�q�B���n�J��џrŠj]ؒ�k�g�r����*��ﶡڶ1��+\�@�����*�V��.A��f(E����f�BB�DA�{i	��f(	�zh�A�繾���̟9��^{����O��wt��И*�wT~���?%)ģ�<��m����o�&s�_p�:w��"���)����Uq�|��'�;����Lm;�ģg}��g�t������(��3�+�P̞����9IX�8���t�![��r���/BK���U̥B�0�!�����/�_�k���l�zVZ����=�Ŗ�NV�I퍊\Nò���H�,�;>{�(�������\�����˜S�?|9���ч���lR��lz|��TWd�'���SF��E��$�N�`��w�X�ٲ��h�ڼ������[G�o�U-���	���p����b&��	��������է��X���@YC86��o9�=rټV{�'%�Е���Gw��'V-ƃO%wU�z�c$�~��?Ir�4��>����<��&�:T� n��&�Y��~h�'m�ѡ�_����8n*7����B�ê����2w�E�J�3?���e6m��Ӈ��f�N�X��ֹ��~�a�p�:��%�<�%]�D2��gb�2���I�(�[�O�o-A�m���=������ܻ�2�2���UR��?��{�I�<b]f�43+|��2�@h	�q˽��uV�!k����2���G�+N�{i�I��s�w8	:T�Z�#���r@q4y�u+���Ƅߵ>�SWu��䌜�n����t�I�;�vX�U+�ǂv�q-�agQ�L9|O�c���_ͱ�t��Q��)����F�-1��U�ڴ<�s�$T^SO1�K���&Fu��&��6��|W�}�P2�D9{V��,�f���߇w�2�2�C*�p׳^w%���,���P sUw�.);���)j�4~�t��T@Xk���Fm��0�b�����S��q�3.�ذ�M䧅�%1���"���eݾ
�T�籇���n��_��ȚR!$h��xD�lZX�	t��7L�oӬ�:�>����U��������@�՚�x�=o����ۀA�f�ӌ��C,FZ�Le��?��["\V'��	��uS�3ȔI�RS����I�ՑO	}����ɑ���³�0����C�r�%C�Ig�-[p�˵��O��)�_����U�uݪ%��
��HT�Y96|g���Ǖl�����XR%���QhA�gL�T�$D�@T�MۍȊ���=DM6�~2���/�X�Y`ʊ��	��!w)΢�[1�u��NU��I/6_�қITY׈�8��ÚT��N�ea�u�ę/�����̀��$�sF���5�)���T6���w���#������z�z<R��#�*J��靸�ǜ�����|;�6��L�_Z�YL��@26̔կw��������S{(s�žT]��{���>�j���d��D�������/�u���p{+�)��w��jn���P�^���V�������<�M����
� ���]bskQ�4Ro����u��Y��A�aj���л�5�]∇�{�FB�+1_��pp�c�c'/,�+�o	&u��^���Yʻ@=��F0<Et��J��YYI��|c��S]K3o�:��	|��֎
���ur��X�9�D0�ԃ�K���-�/q���,-�A�z�6HA
�I ����$8K�� n�n�rleI��}��_,k��U��J"�6�х>��S�a��?�)��B=�J�zVNY��cf��5��v��3�b?��Cc#ļ0HqI��L�Y�vE�N����3���ݗR��uɁ�?j&��Q]T��,^�r���v|%�\�>�о�!z���7�*�%n�gn��|�'�J(�ɛ#2���#k�{i��$p�\�ȅ���X�@�T'����l��O霈��YڰJ)��H�bOBU|��^���d�<S�vZ�K �m�q�A��u�`����C{�s^��H���N".o���b�	���+y>2o!�٦��~C���Hl��K��:;�LU�Y�[��yg�귎�;DsPM�n��D���#/��/��ۍ��=.�����?�)3S�7�3I�����k�j�xP��W�}��i�;�#��{�]�D���+�Y$���6�GWa�z���
+�����z�Ё��߹ߊ�X���_�ˌ�����f��UT҉5;T��f?RmJi�kx��/@d�r��Z�"r�z�)�U�Q�o���M_O�޲�Gk��8�^���q�C��.`oeŗ	�R3A�%'̫��d�IU�����[���ɚ���S�A�9l1*÷�Ҋ8ف�{tf���*���n���q~�:k���

H���4�&i�4�׭�~�5��-�z���.���60�'������w�45B�
�n��C{	 ���������So8��n���e9��������O�5և�ǣ3ر��7�����[��	��K���;�*�q5	�\z�j
�3��R�8��Wh]DzM�����"���8Lc�����@U����^,C:,8���$��N��*)G�j�.�4|v� �N-?�r��5r��l���[M@�E�'{[��ɾ�U�@�G��8����E���G��8���G��YQQ�� ܛB
M�/�d��V
���=d�%?
jYw|AQ�->�R��ƏU����^�Y��g|��Σx܌Zޭ�и�؟+�t@�K������m�Z|�]�
��H)����:�\�B��������v�]\k�����iʆ���-�:.kT��YX�m��*��0g���$M����2�T+��S^�&���w@��L���K9��bV��w_�j�AthH��
��uȨ/?S�S�������Ϭo�ǃsk��(�1�-�X�:�p�4/��9�<?�R�j�AD����`yS,˘}���8:����%��>���(�#�fV��).�������nN�8-D�$܏O��H����+���E4��>"�5���0V�|�r����/ٲֹ��+���a�IE98#Ut]�f�2ܣ,�ʻ��ړ)����5����0�����`*2_�`7C�]m<e���F�µ��}�p� T�y�O�1U��:ݑp?�[�_e���{�շ��M�}m<"�NG�>��I��6\�c��� �
�]r� ��e�����iE�Ʀ�gJUiEnj��R��0?��  ��ef������jK���I��#$������p� ;��X~&@8˜�1#J�fMÀȱ�V�t��	��(g�XY#����7�g�E�9ծֲ�Ψ&�����=�u̲��SNK��Y��Eɸ���R���+��M�c�z�,}�zY�W�Cy->�l�Ya��AK��"O�̦8U���X�>�Qm�%�m�<� �x�?H�]f�3O ��d��hr� Ex�]��*��Ƃr�Q�۹+ �K1�'��&=K&6���l�O!����������]��]��s't�<\�5���q�^EXҖ�)���<⧼ �	T���~��.: �q�I����S�C�ڊ�_Ǽ��ʆ�ѓ7�ZsT�'�.�3	��	�&E�rE�o�nfPl��5�c��uVz��(kR�W�t��ɡm�qIx|�q	�������=x����5D�~ sAiU��b����Q��JC��J�[f�ZAx���|�	�+$l�dW�/f�����!.��5��ˎ�~�W�0����6[/>�]�{d�7]Q}l�ܺ�1����{��Զ�Z�ﭻZ9�yAݾ�F-0������!���:����t�oZ8����������Fi4L��~��:a���Jv/�Ip��UEҌ��;�7kگ�B��m�=mV����Z����k36��W�	oXg��i��?��%�b�
�i�bf�t�1h�C����ަ�uܳ�������ț� ?ǲzV�o\eǩ���ٛ䀠��:~~�����k�&=8B���E�ԩ�=K�SwUJ{��7
=:�������5M���I˛ym~�w���f
;̬W�l��}8$-Z����N=����?秘�Y����V���_'j��C��8����ZM5���#}��z��oa�r�W<�r3<<�����eHxp�8�>:�o����z�^F�7��E��}�2bbb[����V�����m��~��G�}�":�^��թ�杪��"HZ�4V�4��'>����n;L����:����!55�]�M����:eK�szr��;��B��a�a�m�O�@HC�]��0��b�����O��4��L�)I�[k�;����qDh��pD�Tk�_�ߴ�J�,ڊ%������rd�{��pf���z�
"��5�&o �AS�/bߘ=㖙b~���bs�`�6w�i;fi����(���߽u0+xC��
}��Q�a�R�J84+��A��.<���z1��c�ώ�>��Q�x�<|�a^#�h��6�w,���y��@#��yF,~�<�QʿL]�?a��c�;и71���"�20Z�K ł/�q��,}�W���Xh�{��?	�*(X�Zp��so��#wN���ޤk�)\�!$inl|ӝ�o�����`�ֳ@/��y�>�q�'�������݈�O|���	�4�<�X�A�u	p�"���O�x���k��1 �)#0�{��a$�z���e�U���D�,)ÿ�2z������)Q���7�"�?����f��\���>�ٞ�^�sQY�>���ӕk�]���R[M�a��WNT1��$0�U/qF��8ٰ�.��b�HA�A��_�jVv���<n,czP/µ�����(K�s�/�����V'�P�nڋ|��}<F֞�ڵ���og�P޶K�g$Yo����6,.U�w����	h�pcf�ψ��,���I�b�_�>m����ʻg�PC3O����7�{,c'c/�MbSa���ċ6��{c���Ɔ�Y+%�"�i}iR�X�z[yŻƟ���a>��)�iD���9�^w�[�8QIg�ŧ'F��Ws��Y��],�bB�cHF��b��/���|M��g�S�Svs��M:n&* �7��t˱��fS|���~LQtho�Y`Q$!����a�2YN��'�(v/"]-��]�0nW���_��b�@ب�����*��"�zNuU�մ�g`��:6�7���'U%����م~�zP�[voG�x�l�_�U��R3=��� '�ki�1%�Y����:rꋾ'��}8�	ˊ;��шE���Pس?���7��3x���I���>���y���tQ��"��K� ~�.1��4���5J���?��³����J�`$lvil���"B�ǳ�Om�-b��ʁ�ZIY���y���Vn�����i��;o;��=�z�t��u�d;6�I�-zj����M�݁�@�7�<A�^����o�E�U��baY���#_Bmj}S�R���u��Z6����7NW���z���b2k��B^M�����_�k�PP�A�Db|�19�A\�E��J�n�Ix�W4�/>C~�-	9�_�Jɔ�X�B�MѸ�=+�����t�u�������z���4�-�{p�ML���G�,'Ye����[��K��|�$�={Z��%�ny��hY����R2?K\r@�7U�����E��ƐE���
�t|q�����p���O�*z���0��z�Tt���@X��%��'rߤ;��[��5�y���^���=������l3�W���5�̓_�8�w6��/C$�yE����;k,BX��e�|��0�X<�T|�>�?�	�x��I�Q%���7j8���|�m��K��5������c��WG;VY�AIͥ��j�Lש�q��,3iM�SA�a^#��R�UJ_�4Q���7��K�b\�Oc���>L�����g���'(�H5f���W�)d�߄�w�ȵ��7�Z��B������f��0��`4�ܕ������;�([U�=��<�1����l���3]���g{�5�F�i���oթ���g<N��X��P�%���.���A��b��hвq�,���?��Ԭw�j���n5�ԑ�+�\�>?����|�u�t�J����U��G}.�N� `yZ��O�Q��~S�}�g��dF��`�4�Eg��Z��Iډ,�,�U*� ͫ<5X�A4P��>|) �|���>/����R~d�eDC��@ͬ{(�
�>�ZT�.º֞��-.��ao�m@3�����0��X�@w�7Ҭ���`���5:�y�N^"f̼�V���Xȹ���p�[���x������΋-!#wa�e}���]�>�z�iÐ�N�n��1�t��"%��~��u�wb�̫���r��5�7�Z���Q(����%CCjum�����Z�h9	��AGR�Whp��u�2�8B|γb�o<���,��7y�0�� �a 4�d')�;�u�J�����r�[���8�v�Ƙ�l&���=L�R��!#Ѡ��O���Gm�ҺN�����%L��Z�RoYo��r�\����(U��kk���Q0��=4Vv��D�U��0/�!RN>3NJY�h�2-]���i�����W��0V�<�a����7j5��&"��R��j�)��s6��=��~{9����8R�A���e�ݘ��Le�N���0�C��&D4۟:���e�D�ay��Dk)(�X�gj*�Vz�ů�f�t(/~#8j��C�'�E	)��2�M+�ҭ��x��z������֣;�����*�H�V�J���4�~ 渘����w��9����R��h���Z�F��&,cdc;
��Pl��2��\H=�#��i�A�`~/ ��s�|����Se=w������v����[�J�.�č�}HI�tKj��Z����2I�p��ZvW�TN]�n�Ā����/�̛9m�؉D�XՔL9�<�o�0���:uN�}�U7�i���',Pl�_MM,SU��)Z����y@��\��/����"y�-���(���y�P�~́yu� �R<�ԀO@�u�a9沦#��Td>��{ݳST�8����>/�S/,�>ƫ�"���٘!�4��
��4���p��>En�bP�B,�у=��g|�*�9ۋ��&��/�B:����:m|�C2d���l��i9؍��	G���_�<���b��փ����1���i�P��%�ǥs��;�q�M��*�K�4�5�֒ͺZ�Cɻ�}�����Y=u��8{g4�)��~�e�mVf�g��Ҙ�Uf�(��}h�^R)�����M&G�$��m����=�ܨ�{��bT�O&�w���t�ޫ���!��÷3[�X9����E� 2��z4�s���.7��4?o��+o&�7*�8dF��+c?��I�}���A.u��p���������{�?8�È���疠?�7��f{<W���9�5��*b�i�WQ�������o�!K�V����`��
x����G0������vd���楶b"J��]���J26�A92½���C7����n6�d6Ms��)@ZK$C�ᕈ^��5�w"γi��ח�1x7_ '�ZOa�y�}+3�!���7v��r�	���=�$e���e}l=$�?�Y�����\�=��l���zf_��*b-�6�Q��q�Ѻ�n�9�2b���Lc����礓
W�F�c�$�9l�
u|�.��]R{��q|W"/)���}���.T	ٳ��#�T\��1x�4='��w�AG:{'RW-Z@�v +�j5����x���2��l��e��Y�; �bnrHu�Uv���i�
��<v;;;s���18�M2;�[�{|��2%/�U�C���-�
H��f�.�M�'.8WE�uQ7��o��2C9��gIm�~|kj�԰I�hg�75�Yyxŗ�c�*g�nw��}�9m���Y����83OXG��008� �푴A���~PY�C=�u�����_�#5�yp�}�I�� ��w ��O{�����r�_��!�hʯ�l�-����qoڪHp�"zt�̴�6Mr�e�D���2J�I�	�N����j?*���� (����a��?/�d�$�3g�02�Z��b��?��mJq�}����^����#��c2��P�h�u�qq����oE��a���W"j���ǑI��-U��K�[��O��	�ond�O�&29F	�w'ܴ
�%#�+�^���ӜIi��Ȟg�~�f	��M�T�~뗩��{ g�I>�@-�B�X�߀���o�ا�븿�n?�0L`����yϠ!���q�,P될q���3Q �����F�p߈қdK��.xNA���U�aY�Ӊ�7��w�䯫C�����i
��� u&!+�1�i�F��k�Mv �[�:�IbTT������$���ƧjV%����s��aJ��0ޢ��T��"�X�J����]�k���ˑ��b��+��=j-�,;m3���-#��[�*BS�4E�L��J�n=?��p�l�����o�����p�^d�j��
ӏ�b+kk>��'9�;�
8T	��~���2�-wT���46�p�y��4�ֆa�U�6>Rs� ��y�L���F�K��}TF�c��*��$4�_���s5m]���R��c
�>�E��: �J!�:���t�2���4�.�[��mlX�.�giߞ=-G1���6�-�U�Zco/K�+�o2H%2d���u���}����eӥ�i�%���e�H�U�<m�Ư��S��ъJ�f�ce^�?��8��t^��p��0���n$�}`ո�ʣ�T�5 Bd��:�ף���
�{7y�i'��@u��)��X�	�Z�u{�й���F�ۆ����ޡ�̿6�1X�k�KH�JH�N]�<VId~�
�
�2VϾ[�h�?��g򑼅�{yF�L��D�'d`iŀ[M�n&G�#k)�e�K������f�/��=�=�d���3��>�%X����
~f晋]�ӊҲGS����~A�H���<1�I� A����������BDB��k��%*���]Լ�[7�Q��X�i ��whi�g������g�0�C���"��]�f���2���*>ˇߌ�y��.I�T��f,�U����Oߎ�Z�W1�06�\n(e��셔R��du��1N�嶫���h���G}��X��w��q�����~�l��� {���l�5[��ہDv�Az�OnZ�f���;��W�
D���ׯ�"�2O��)~*��3�U@���|����KK��I��È��
lʫ� ��	�S��h�+�Q�X�h���$!A��&� 0��3��vY���=rN:����u+:*wY�����Q�~�I�KxE�EdݑN�ܯ���>!������#�+�q����&��oԹ�T/��1�w�����_�Ft�D^����2Y�����6�9j����%hRH	Rތh��A�/�`ۛ�ra��ZG�����=г��ExM<�y��=\����؇��%�$��w�N��d�u���ۄ{PN��b���+����Ne���
�x�{��r����}]���Ayd��?�sh�������L�\1�yL��[Sz�G��&=`���׸t,;��fɄ-�M���۩<�K�^�#Veggۉ����o��#��u��S�S�B���� 0|�W�#�ۗ���~�&�+*$��ZLj9�:4�8�!G�T�S��7ٟmB&�L
�Ǆ��8���M���RE����}]�R�lW�߮<+>"�>�yX�yd!��X���
?�c�������s�e�R��rX��Q�s��9��3w��)�E&�aQqp?���� �5#omMG4���E+���%�?D��x&0}M�d?�h6G9��
�I��%'2�j$0aHj����W�t�ϓ��0���:!|���Ԕ*Y��g>h5?�̦���Ŧ'
�:Q�εg'�"�_�,0�[�@��\>\v=�,ϑcǅ@�chB��a&X	���O�]>Թ�QK˸*V�c)Z{4�-ځ�?b�m����6���tE�BD$)�_
�hmOMi�H�1���7^�+@��Ƣ���'+yv[���$�_^�&Z���n�ݑ;/B%`�%��}��UZ��ZN��k��k�Є!k�u������Ac�9�z;EÚXD]� �}�͢����Ï����GD>��]<���-f���m(�-�)o��?��t�����C���|�34O}K23^��D�;&b�v���T��E�M�����Nf��D"�K�o�-�;k���F5C^��蠲N�2�^�8�U�H6�f�����y0K���ڰ
/թMG܁�z��&����[���d[����)����.�6Vb���AxG��YKl�W~��wH5 6��h�D�L��jV>=��( ,�z��o�MR�`i�Y�[����ad��j�HS���M2b��[�xg����Y����3)F�t����eN�ZK�%�~ �w3v�eC��?�ʞ��&�\^O؇�x�r�:X��XK��u��a���3������[ʀ �jM��K�q��F+D����|iAQn㡲�ڽw�����ɓ#�1�/Mg�O<�;Ӟ��36�c���#�߻~��_��k�s�y�ʶ7~��L��u�w�T���Tt���s��%:�Q�M=��=���Ԏ�Q�H�9��� �'�\Ȣ���Q�p@���� �_o�H�n�/"b����v��*�5��>�f��S�k�V��y�:�W-�R��_�AY��qxxxZ�(�Q�Ry�������A^�����
G�[����73�3�#���7���N�5!j�z�r�󧟣�\ K�^�eo,ӼsЙ����3R�|j��j> �uW����N�`r�+s�*�Pur���#��*1�h�]��+ a;@ݝ����7�8��h�!d'�E�@\���l���On`��^>��K�42D�z��=T 3���l·">,&�Z����&b����a�#���o��J�ť�d�\J2Uq�f��jL��3-���Xz�Q��2�[��<�C�Y����Σ�*z����ۓJ11~/1�ꌛ�r�Z� Ֆhf��*4e�h�P��Ɓu�/��C�f�B�?��o���Z|� �m��M�^��)�7ɗWuum��~9���˻��֡��vl�<l[��$�S�e�+ü4�z�ś2颕�^l�.� �U�
*C��g�9:��jh��yB_��;(����7�CP��M(s*��;� �5���L`}ZќM��|��[��4�
�����* ����_�i���/�ͯ�ٺ�a��o�~[g�(�dP��Ö��m���6�0���xc��_e�Z���|��ј��C��X�4�FJƄ�:I���S[�\�z�˝�_�����}UqAՇTtF�V�l�AF�;(V���4�uǒWP�b&�&ɡ��c�V�4����{�� m3H�VW��*�ÂR�z���VX��� ��k��׊&=�"�|4r��ׇӏ:���3�$,�N�@���#e�����W��y�s������Ҝ���q�0��<%epz���+�߈]D�\�OqU�X��3��a�QE>�+���ER}�J��9���R��B��G����c0���b|�GqV�z��]�X.�0��8��Z���U�1�o��+�˃�i��ʷ��@�����Y�㖐�o,ٰ�_"����<ǣ���*�M���,��i��	EqQ�H@WH����{X��ƓO����P�U�uum֡�ݝw� *+I��9Ľ/��A���I���i��s�v�G����Ɇ���_y���.�x�9t��\�#BV�|I��R2�������!/�7�j��G����ΠoL���������8�:�%�4 ���LH�۴��SDM,���+5ni�-��8����/(A��5����,f�3ʤ�ʪ�v�����p-��喱Yl�?��X�C�;sV���N������l�] \���&أ {(��s��j�Z�ϴYzݠ���CV�D`.�Ğ��'��8��}������$�c+�F���~�����~סwU�F�w�iC��\>Eq Qד�9+��}Yh%3�/�U��^Y�Pr'�������c��:�;*�\�0n��@�d�'�t���++b}]�?J���[���j��(YԄ���k[�w���E���%H����I~��/�������ͺ숙~�d�﨏��L�d�%6%��/�*d1'u.9�|�aFS�����)��YA����d�? ���>W�)E����t��x�~?ow���#ɳ�VÊa�`��B�������>��6�9$I;������?�뮭�����Le%wq`J�~�d�E�v�-��JN>0>�Y�W�r�[��X�~O����"����l�5#G�83k�{
�Ӣܛf�%L�?q�|����~���)<T�N�J��PG��Ki3�����!�/� �[���D3ؖ#�}HL�3�᛽X�����Q[�n_|��O��!�>�v�9�ilSb�����@��y�-fI�33l�wG�;�j�����s�?6��;�bV1��#���y(ՇRfU+LJ'^"�B��vk������B�	�$x1�uy(j�`����nce�m���a�Cf��l�ڿ���2vӠ��Zm7Z��H_qZ�P���د���3$�v.���.�SU����;�ĐrD$}cٷ&P���y*x�Lw!��rlHL��a�8��>�tM;V��͍��D��W�c'ݙ�<)�>N�jk*���%G�8�4��wR��w	l!���`dR�AW��$ʿ-&��f����2B�������o��.�����_uG���o`YC�M5=��$�z�H�.bS�sC��e��/�Ї�Q��+��+�wD����l�k����'0��C���\!��P�)v�{Һ��u�S���,�>F���}�B�� 륧k�$B +�-E������>�j�A����>Þ��a[~�����ǅ�����]s��~�5�3�UpY�xw�6�	M]o>rh�kV���:w����pu�l���Hxe"oؗe1%��P'U~��4� �
��g*�&���c��3�b%`O3��'��y~��TOl5{3���wm�s񀟯$d��*���6��*��Dx@UW�*�P}�5<�)[��1����Ow��u�]�LH8ӝ��!j�%�_��ܗ�2�`՝���tԀiv]�C6%d�K�Շ�H��zt�w���Q����7�e^�.^[\d�пEZ5�<j�����IV)�ʊ�����$�<D�-��_lB��/3{��"�0��bp"ry2+��A'���K\� �jNy��:�H+:��蔳EQ�[���T��q�n1s��rx3�\��W���o���R3`��^�~r�O��5�j�H���Wj��w_����?t{0Jh�A��+Xh��L��`1}j	��5z���'�A���#�c�d*� 'A�\�f���#b���JKP���Z��9�վ���'Z�^�/.�98�r^md������2�x�.�n�φ�������YG�G�������'�)@9�����/�@)洆�D�)*�CB<��O�d��H���	�5��ʀR'|��uZ�%^q�W��N�X��n�ⅨXt/Cg�bݢVp�[Y^t�+m�A U����1MF��&O�3��-R��Ӽt7����d�4��aZ]���U�Ȧ�B�c���{�Veo�a�H��J\ȣ����oRk��s%e�[qi�%|'�;+�3_rX�
"vGNW���|��7&%���ߤ��k=11����m��:#�������?ox�+8�/}�c�}ߒ�튉����\�*��A힇چ�s�033HW�?�%F�UZ�k��R2�t����CC�({e������e	 �}�s�Gwj�S�f<�ƭ�$~��O��]��J���B�"�ɷW�O�ϮAM��i"�sv���"�yS,��=r��s,�L{�5,*� �p�  �L^8�ԓ���,B����*_�7�4��/�3����42M|���8�8'�+9�6�%�λ�/�z�k`�7���]��J;|�S�5���A�m���������u��iR��,P�&��zR*�%"���B�kfjI[����c�'����B���<A�T�°��${ǩ#s��ܞG���3�U����1w�L�x�\��B5"�mV/G�]^�z�2����o��|�g�����si����?��z^{�B�%z��]5�+��/�iXZ�T4H&�ht���ڣ |�Y��x���,���0PG;���0r��i��2�^��l��x�Jv+�O��N)����T���<��FP`��%�o�!��&���Am��ky�%�߻l+�8H�l�
�/��Uz@c,�ư5!�8���52ɣ�����UEX��ӷ9�˭�,��M p~�4i+tకU�-]#�l)�GYQG7���Uo�>}Q 5��M9�B<�J�0�d�w�8��Ȩp4�:`x�:��j#���^�A�5��Zxe�IďjM��s�ƹ�=����x�1C���"j��dk�oӆ�j��S�������^����l?��-5B�yW����KG�5)R��r�`��XxAԜ���	�����wrN? ��YI2�����L3[�r6��V�u�?^��A�a-���R)i{2pS���f���~D�~%���
��(?V�s���wS+�����_vU���c���T.)W�q��`
)��oը���ϯA��s|�Dt
AU����%@E�J�,���U�^��39�t�HT����v��<��<؝>TD��-輄�m}��Lu=+�]�l��T�
�ɡL$�u)#EZ֎*&a ��� ���?��&�'��X���D���g�j�%��o��	_%J����D667� �� �];�=��ڜ
����/���E��VÞ�y��i���~��	�u��MлFz����W�4O�.O���eӬJ���9��b{�/hxfh��)����wp =s��c��Q���n�v�a'��)!L!����ϗ�,���Pwi��6_�dD�)�5 ?����p�X��b�R��|���!q3`o�ޅ����� ��]P������ya�X�p ������SI����u)|�c_�(�7�#������O���
��zz��(���P5(�X1�.�bU$¡'T�-�;�FE2ь�NM�$���>�UV�w"��[<s}���d�=��rW����޽�Ks��V��D��{ܕ{7�h" �ń���{%���^�r�i��>���0�Hr�JM�(�[4�\<��'�-=���=�&��h��l��aLs"���?�k��~1 z����m�*l�a1���?�醙=���n�N[�k�Y�e�"�x�U2~���O������A,��G���x;��nU�����Z��˝�峒��)�e%�l1Zܛ�Ȁ���i~7I�T�2�z7"�-� ���C�
��_蕼_�����0hU��jv�� �������g�t�Ǥ#P��󿷋(dǌ�\��rU_�P�J:�qD����'�<��H�U���%�]�TUN�`='�T� �=��0�
�K���c��6e��Q��'�N�+�J�!�c~����/�1�rd،p^���"��&�i��pcƐ�ꧡ���K􈾟=��{�@�`�Z���N��,x��������p��%������̻wr��ܹZQ����� �f��aU�K��jcL3@�̟, �U0��L�k���>�YĆgTH�w����*K�p�n�=�4$E��P�㷺l[UxFtlp 8WA���Y��-��g<e��yNd����$k��Y�ӈ𻆉�(��͡|�����v���"��ѽf������
���'ݖ[�'�I/�oз��wV�s�0��u�k�ul=Z�r�u̒���	�K�O������{�z������m޻�,���j^/���3�<�}�Y�OC�ugm�A*D3�8����q�c*kz�Я��V��r���lR�{�k���/�sa�+6�t��8ӎ���ƔR=o���o�)�0W'��q�!��<�ז�-�8�,�����;�|��P�l�g��K�❱�1]h�4ԻP�yK����>�[��/3�������Mw��I�l�D�>s������mp�޳�59������r]5uuKGG�TU���|>T�U2��ꢟ>�Ud�2Φ�����Z��l�
=�K��T�4�Э�p���x8T�w�b�&���D�\��4#B]8�Ӧ%��y�A�s5.i�n&�>mU'���5��j���'ٓ>[���j��C�{\�d���a�����#��N^AW�nvv�:��Ƥ�ώp�Ʉ�s�V\�櫛�\ѹ�w�[���_s;���Ͷ�����!��N��W�P��eb H��R�K�dd�.�T�ȕ6�Ȗjk���ՙr]z���;u��r�	�&`6��s���ɔ+Gz9?�oc���L�h6��5�W�iu���1�t�Q�:2��'��:s��>��a���r+��9�OBU�n�t��m�,����9[^.�5X��e"I���)5�;��[s=b�g�\�M��L`'��ʚ�bᜂ�~�c'-��Q#M���Cb��el���?G-y�a�E��������'^����QQv�ޤtJ���t# ) � !�"%� Ҩt
HH#��J#��H3C����u�\�,������>g����~�����w��qț����Q;����kO����[�$oo�������K���"�|K�= �$}�52%�nw���;����eec���UϜ�0�;���0�7۵�����A�����,��MT��~��"MJ�Ŵ�ʮ���S7Ѯ��9�˲)Ͽ�l"���#�:����aò�sM��fb�����ô����Pl>~��S8���63H���	������6/�:��S{v�EJZ�.o,Yf��i�#`'��|�QG$J�J�'Xc��\��d5��#���) ��K����Ff>��}� �Jz�7�X3�Gk9[�"_س�E>f��Ń����]f��𴴴\dZ�Vs܏���n>~l��,��a� ���ii���%��@��̖Z���xD�R����*"f�r�b}�-R�8��}��Q�(s�!9�)�۽��ז�8
�Ƣ��.�E��A�������>�2-H`-G�tF��($���w�|Q�tGw��+a�S޳�P˭NP������hL���Ԣ�� ��Ym�Qm4�	&))��������e�qV������#���^���с�Ч �gnVu7��ƫv�O:T)c�Q�n@,��\�fJ�H=<<$A�ÙOC�i���J���g�F���fJ�ah����u&~��x%&_���}d������s�ǣ��e���n�<Z�C�]�<��c�rE��褁��V̧�Q���pU�i��3ㅯ�$��4t�G��� /��uyN��eL�f���6"�OMuup�f�c�K��(d��<OcZ�Dٿt�44;�ҠW�/)�̄3o��T����T�^W��2q���Z�tKv��6�՗s��f}b�@i~pr�����rfaNk�]�f ��2j7ˢ�C|n�+�J%�/�4�e"�+4��-�%Pn�ʆ��7���^;T�jO�trf!_7��q��I�s`�m���ULrQ���|j�Z?F�+�0�-����+��u���[�'�9���?g�m`X�O~���z�9�w����܁9]�����s�*Sh��U���|�s�D6�)1��b�[+��>Z��b7��k5����X�9��o��k�eh���0��Pk�?��D&ઑ�$��ۡ�!�S�mmquuO<�lV��D"�ūm��UU�Oͧ� |Y�#��o�t]�F�ܛ����L���_ m����o��j1F<���+yLo��Jj�'h�_��ԧ����3z��7H�$�F?�]����^<�D=+s��'l��w��(¶S ��"��5��ȡOG$���x�@ȯ`�����>�%_��)O��c��4k�D���I�(U>�
잕�;���X��,�N˿�Z�)&��cҍY?�.P�g+���Cͻ���d����_SO/|��n�c?�tuu��^����>h6���Ԅ��ޡ��u>�WCS3��sn�=�A�Y�Q�^�-^�3vK�����@�Ufʂil�3;�����9�^V�:�N��B�}8��YT>i'��怲��A�!E�x�-&F2�f02�e�/x�
<�7��c�#���u�1�����;���>�Pbt=� �� zSXD�
�1�/��X����67�.\������nF��(��<��HWF��]��ߠ{�3a��@� 􀞞��x�bjj���9�/�y��@�nY�g�St�C�`�@jNN_��4:gL��莎�]W�*L�ြħ_>�)��`~�jÇx�9�����_S��wV�J��d�AZ7��ٞ�*���~���9��b��Kk<���q��M;��(�b��%4Z+�mt��ay�ƶ�gE�������5�N<#r*@�T��.�\1*hZ�L��UiZ>�DYZ.E�l� nĽ��M[�oib�e�ep�,�%�7��[�����M���d|q��_  <<L�-�Z��@7&��� +,Je��g367ﻸ��%�>n����Y�' iMZ|(6GrPp��GF�M"����t��]��h�g����HI���h���:Z#hF����A�G,hAY��/ "�(����f���lŵ�g����׋1�x�,��p^�%�E" ޘ{h_V�;П~k��SnI�F�O��A桄 q�v�n�+8�nL���|�飈�>��w�]u虁�3������66��L�y˞݀&605���q�����z=�1l�A>B��T��1]a�Un��z��O��F�-���#�S6Dx�����W*OВ�2YŃuٖ!b3V5*;�H�}��X?��4�����~�F�ֺ�8d�����}�S��c�ZksZ���<'ǳ.j�l'��˝�J�S���������>�r{��c������^*��r�g��ֺO�6���}"]A���3O���D�f�̓�`�吻^+}�;Nd#:Q!~�h^mF�o{J�k`h�17��I�#]c�/}�X�G)����)��?��]Ox*���x�+�C)��{{{��2�T�"�U�b�S��`�Xꅗ��\̧�;MJ�j�=�o�}>��J�1�_��{�>��*�<pd�,�e���a叝��|��$~U˿���� 	~�����b������`��қpo��^�B��%T��`�=�!"��Oaܟ%��9���Qr�|ի���ᡈ��>�7��m %hii���-'-����X��ֲ$i��o�f�rC�u�K���Zo,}�����|c��t���� ��F��CEQ�FɽI���ū����l��?�y�Z;-CstAA��ј��7Y�Zw�Ozo@��ˣ��C�J�ls~N�ƚ55�2��~��C�rys����;z���@�O�(�ڐ�� r���đ�;�E�9��Z��&i�o��Cȿ������#\gD��a���������r���wAe�k?sO�M���F���1A�t����,�JMH���Nhe���/%��Á�����ttt��<�4n'V�����Gypx8o�é�M��+�N\�z�<6C�J{,����N�A�rV�
�ɓ7y7�Ƙ8	>��*��x/SD����Ҩ�9����$Zܺ���AOi�$����=`�Vf̀Q&E��:7%H^#s���� (X���M�8Qա�;�ڢ����v;��/N����^�&f  �tG����4r�t�����f`b�`j��'���P<����s��t��7s�Е��K�r�I��vO��oZF�LUܲ�c����l$^��_nk�9l�nT,py�:�ȥ{ѝ0����\+ڨ�
p�n�~|i ��hG�e��Q��y�=��WeQ�L���g���۳?~J��}�nnL)��w]�����%�������K��P�w~/�Q�E�cZ�R5��+����^6�{�ō���~h�������$Wpct����Oԛ�����f �	O�1ȀO���� ����INIA� �D7����(n�ۘ�r`�%������H�p��Wfw����i3�+i[�7V8K���F��_�џr����h=�v���	t�l	8�ep�K��COXxE�O�G��m�;a=�@2��F���uV% �~�[��%ߗ>���c=�`VL�2���)���:��R@�A���%�γI��P�/�^>MA�#����m�*����p�V/�}ח(�?�9ܢ�����H��@�q�L)/B��cJ��0t至�}��S���w�s��v�PN��p�q�*X���=t�2�8K��l�Y��H��|���^�^D=�gߓ�����[w�ۥ:��";e���Z�k��j���K��5�z�T�f���N2~gBcsJj]�Oh� T)M�����_pnb\���-ݭ��L��y9�_̅DD��RgȖ��(U�I��9��?�)#7�aNh�$���Q'j)p����Kv{7���R4�E0�[h��<?����:�Y	�u=���voڃ�`�E��������^��MlΣ�~�]��}BV����"��~#�I��%�U��6E�#�s;�q52ɳ���yG��`E�N�����I3.��Rh��8����ӿ��j�u�B���G�<[˷,�z�<���b�;ńz�6����ɴ��2f�徴�ѐ����L�&	���M�s�g(�����bk4��ň�����m����h9aǉ`T��bum^�*���XX�2jE��C�,j�S}8x�z��NAꣃ��W+�?:ۦCͱcIb[M[D[�����&5��j^����|�Y����7���	����򙥚�������b����b+���?���i�d�>��������>\����*��4����1��/ƃ��]s����\�1�����O� 	neoO@DDtv
sAF�_a���S���ښ߲�����Kk ���םD���_O�]��kQcHB�������o��\�>�]�uchb�6v9�r�=���`gh;lv!�Ȟ�i���������.�M�,!M��j$�"��;��l��j��^m�r�v��W�/뙮�����S<i�@���O:9�ϾȪ���Y��6?�9Io��u<ʬ4;���<��I����� �c'��ߗ%���o�<�n�71�ۥ53%���A��pX���ry��xԫ�]���4	{,]W���'�ª6�L��ʼ�
�^�����5���0�@]�87���Ah�ǁHP��5���M:���y�(�v�m(_�.��I-���gE��6�2���w����MЋ��vpg�>4)}����i�MK�S��fg�ox�+��kvN���>�D�ܙ���E��:�����3�U����w|p�S�l�8�7,��\��)�uF�?)DHOQ��N��((���oֱ !��	� ��l�To*���$�ഽ��v��7��-���=Q��Z1�����P��}ޞ���$�Dm�ry���8n�\�Ϣ?��%���{�������Sy��"��*��Ȍ9l�%>=�t�<c ���\ox��:�������S�r+ƪ�>,�zB���g�.G�ss}yvs��4����O�a�ێ6l������4�z�T��>48��oӢ/�옂�`�~��<yA���`�mgC5�;! %!	h����X�G���}�� &G������������e.6lm(-��dI�������^�0��c����uO����tbYe%��.�ٿY�u�N JK���f{d&��!ٹ?A�Tvd{X�_f�M�������/��6��cjhW�||#�)#���`o��-����V3"�55��)���hU�Ԩ�fF�cnݐ�MG�Ю����V�ǩ���?>�=�yJ���5Ɔ.dd@P'Mz�#/3�s�;�������W���=��3��%	b3QOڭOV|��4�^dț�i�"�q�,�������Ht�1Q�y^�M@]ԏ�����M�IK�E���=�M'<�<�	�~Zi����1�gs�L*��� B~ڍ�d���#QMMM��.����=neee��b�;�+�-��5���OK��Ùە
��W����hB�>CJ�wW��
���-�t3]�	������Q�zf���{LWm���ee��}t��}p��'9^�����@�W���N~��g(Dk�j�]�����]��W-7�,��⻊=Z<�����떖������E~�������#������c�LXO���� 0us����=�~KUU���5`7�I�T�rc����;��y��&���m��w������R ���Xy�G#�(��ió4�A���c���x�f1��Q�tKU�^䞴IVM�7� әL���1�K��ǺW�Y=����wa��G�e�I�ʪ�Q�sjm�vn��:uD����I�O1qh�p30�Y\��)C�! LЮ����x����g����	�o1���n9���Y��� ZP���g����Scs(x����"��-&��-�7�u6�����k�h���G�1�ЈH�,��!����s$_}q�}w�Ҕ*?�����^�zD��+J�������@���O���ݲ;�+}(��\�����!~��!���zB�k�Jp�S�o�L���Qd�U���Z�*���=�S��f����L@�W��4�w�_��-�`�����j��Òq�h-�Ǉ�u3,�{Ⱦ�w��r��q����޾I�AO!�M�Jr�%C�D�?���_�-��� ;<�7��%���NH��=]N�����8x���c���ؤ?fXnoq������Qߚ��gU���L5N��7��\����6A'�Qu��x���9�w��F0]��oZ���:Z�̇�U�D
�T�o�(��w[�gp�@��ΰ��9҇
���#���.�'4w�s2e����=2b�-�^S:Y'��/�Jg��7l.�cuɞ�kP
U���s��N[~�:֏�}������1�T�y$�o���_�l[��f�KZ��ze�6�[	~�Sc;R�4h���@�����L�o�R�p��/�`����eHN��;�ݐ�C<w/eCC�ik��Y.�M�6��,�!�Ŋu�J��ٶ؟���G������~H\t*�_Q���ґ��n�R>��!�h�Od�W����^�\��| 9y'N�����F�Zb��U`�i�(�b�Φ�T�������_��my���&|P`�M�P�K�*v善�yź�er��&��9���}`��z�?�!�XhqĶQ�fc ��Лr=<+��U��
����Ϲ��N-�M�+��-�y��/��}�����ѫi���5It7�(' 
г́W�uF��U�q����#�,��L[����e�%���NP�'֖�.���FKԷ�͋2E��O^���z���XI���T���GL΍�&^���yէ/,A�z����ux�eAv�$����{Ƨ���"�~=)ƱE$�/�� ��|�(2&oo�������y~o$[V�%��2�%��A����[DOI�@��8����j�H� !��C�a$Kn-r��-�t`�.Y+�_��� ��������ȘC�;Nv%@!�o(ۯ�11DEE}.��ai���R7oeV���њ��Y�ou���ߵ�v�����Ԇ����o��-����k�5�Z�F��#�����g�[P��{ň5�u��� �v#Ka��L%������њ������r�痊v�	B�.6h
�WK�Q�`�9�-����8�D	6�|���@���_mH�w��Q��2����ƈ����ux��e�E1���K6 A7+7�skq�f�����)o�._^�1ږb�l�4����AK�z�`���0�rn1Q���r��)J=Օ��l=KM��&m��!��b������	$�.I���QXT�1���w�i���V�j��x��B��rR*�'z.��H�9��U@�`lQՐ!8wKWՔ�$cN�+��'�uƨa��ɝ����m�ݚگ�.H@Į}Ք똚�Cgv��C�㱗g[����f���^�1_S�^{]���dw��5W��_��)���#������[��xv��T�-&7VT�Qlz4�]f�vA�J��{Ԯ�G݀];��<q�u3@����!���U����:Me}����C�B�l�����J�!ᛂl����G!*�(�fe#*��{~��U�(�����Ct����� �HH�k��"a�B33�������0��m���ɼ��Cd�gJ:<�kP[n�����.�!e�y���3�!� �}tg�8F����%*��b�����7�zfO�]�cM�>�-���ϩ:-8a���~���CԦn�1�f�*��z������p'?�ۀ�Ҡ���oNѷ2 >�)�zoQ�;�ēT2"J����|���\^b`��Yf��J����7�5:r������*+��+�F�R�t�_a߬0�`��&��|�!1�3���!�,��n����G�o���V���\�{\`hi�k�q�K�!Ѫ����j��:"j3�BT����cv^�.8�H�ǌ������,���$j���[[���������|<r����Cd��ZE�u뽚�`��/���}'�)�a>��s��v�����O���ؖ���U��ꎠ��z����N����b��_���J��"�J�W����m�)�X~��z��a1,��[|Z��-Z~�P�̿9Y��ߪ�Ř���P]�R��������X�3iV���{3���āWk������o�))uW�X��ࠗDd$:꼠��O̬�u=<U׉u�d��Meϛ�&�H��T�2Ƞ� _�ۉ8�MU��*���#�����M�E>��Zܶ����I�5���G����E"�3��c�]��iJ2�o���2?ӟ�\E��ߦ�q1O�x?Auv=�q�U�dUעd�G��\�r��/����M���5i^9^�ݟ��Q�̖ `mq{s��E�o<d��3ݑ����f~H�� �I�����*�sw���9��$�O�x?Ӛ�;�S���pU0�J�q��j����O@rm�$�J�8/m8�����Q�i�|G;#�L���r�� F&����Tw�Ӝ[|����}��lH��
6'k�\�p9ܷ��U� ��O'��c$N��'��Qc=5�(txS%�A�X�E-��`.}Ukn��-���ڪ�)r�~u��C����ׁ�����ؿ�b��x���>-�����KA�����q��.�+�����)��U1��Sm�q)��;�����4;�\��d�a%�Z�O�hꊒ�֗�Lx8(*�qkQ�R�2aΙ�>n��I��ק���*�r��S�����+Vt�b��� ,0�R�s��b��ѱ;3i���+�'�]B���� �F����?�M�W�E!�~������֜�8���,8+=X�P���L����&=M�j�^�
c��I��d�t�[C<w�H��g�僕��[�z�����x����ߋ�����HI���^�v�7To��#\%������SD>�1�5�hee���*w�Cs������?����d:�ު�W%6M��g~��ڢ޹��9�<�8������W�j^\��)8���G+X�����H"��ܶy��B-��rEz�WL�	�,/6��9�R�rM�_��� X�/�^�:n�j����	��7.j:W��w��`~��f��'��[-��������?���������(+4e�8mgV�~GCm~O+�.T�w���a~�%O���G���ˬ�Rߪ�N����3��̇��z����dy��&�k����I��FF��IŜ�)S����)����.ϵQ0����`��f�ă�����?m�}�S�uj"i݋�����؟`"�'D�5�1�$��<:�^�( E����t�d�����b��b�5f��Mt�������t(�P�=X��)���	6�����T�=S�����إ&�
),|lx}�xs�[m�C8����3���C
�Vf��jU�M��[���`�sm��r��b7�*�>�_�EY^���w�7�nj|�Nl{X���N��i!�ǟ�����s��@Q��F�[�f�`�e��b'��L�P',�LS�R#��)�"�����]{V!d� !���_-��+:cF���u���e:��Ԝ�ِB��s��@���'�f�^��J��ճ8?\G��/�/ ޛ���I)�OX������N�����^x�-��G��(��O��@�X�����ß���f-r�o�`�'��<�+����8���W��Y0���u0WT��%��ή8�f�4>WR�������ä,Kه3�ey��F?&��(�JwB�I<g�Ti#_=��Rt�Tx��v$�'�Q��	&��������P]h�����P=��~���?N��I}�X��5̻���J�f�V,r�l�1B��yx,	-$ ��'d��N�$�y�/n���3l�	�M_�M���,�ݼ�B1�W��'����D�.���p���T�C���>���J!�C�v���S��(�Ɍ��7��w�2��u�5&��Z�!?T	���;Bg� A ����[�(?i��Ӣ)����Z����s�:�	h��0�c��~��&���zc�<ztn�C<zi�����c��h*��3�'���/:x���T؅D'�F��Oʹ���E��^E�,N��*=�F��p��k���^�.2�݁�V³(��oS�ܶ���A1!wi����1�=c��x�j�:�C�Z��x�^��������9a=x����A���X��^7���#g
����0=�	�H^Ϲ���ִ�SN�M"�����G3*�Ot�L���E���!�x��������S�z*�A�bl@��a�-gb(Ѭ8�Lp��ޠi#=��B����_Qe�3���#��,.�`TŃCD:�!�|��(��o3K�W�>\}+���K�G��+���_���B�tO�Y[���������B�Z.�p��o�yƂ�M�����WxC��"���xB�49��W�W��<	mEn�����c9=<�u
bQ�����s󌸼�v��n�%�*���E@�����̋�D���co[
pCX,��=�����=#k@'zeWT�!p�� ��܎3//�y1.��&��Yl��m�Q���oi����ʳ���߰�UN�#����bhi>���_�V�f_���Y�U�t]� e�2�9Li��9P@`�A5V�Y7��Q�����O��W��Ab >)�h{�8|^�g����Q6ч��n��f�lY�Y��IIP����d(�fe��P����W1��3/��y��o��rx���apOQF�{�D�ë̇���Do�����N62\���I����g�kS��ëv^�*3n /T[�1��%�D<IUQ�D<�9��!م�Te{�%�CĽ	`�o����hR(}�B�����&�
���0q`b�×�"��ԃ.����#
�?��/�ݨ4.��"o�B�4���^���2�:�Y�1�|խ�6�B�/�lE�˸�┲|�~D���{�Q� �(����lO�ݙZ���Ns�I���یc����*�~N"�z�=�sj\O6�"���=��l�9����T������s�w�o`aV������ �R9cD�a]��)�n��y�L"d�����&_:�8���h�N@{���Yp�f��ч�l��(�Z6��'��3�:�N���(�Zh�K���A�t�j	 �)edḽJ�X�(���16?�&j�
�n����Ҋf�<.������N]~�\�u�##�`q��61J�܈.��I:|VY�-t�!��c&R/$Ȁ�y���:�'-�<������B�XxF��$^���_,]]�?)�W�w� �e|�l�xӃ���}��	�I��Um4�U�LC����߄�H
��S��D�;�u	ݫ����@:g��[KII���� ������`	���ѭ�����_��U1F��J�0@��)狰��|�E�:e	��Df��v�����������E���]�&�e�mMCj����d]�"�.=�mᘘ ����N-1�YHԛ������vG��w��|�SE]os97���z}m����sP(��f����yU��䫲���>7�H��Y,��6K�6����V�����u\Fi韏��4h2F���C_y��gzD�k��K(R6j9@2�/�����}�A���͵�%����g��XIrb$i��{���u�;9�b�����{%�%\�"���1Z�M�ۊ���� 	��� b�XQ\�Q�/��͐�[��j�H��U_<�e*�����+++�\گ��]c��A��!:�������쏄���O����-�E�bh�.4�8�W�>��m��=���'�����c��L]}�|�_�"�<o�/�8��J5���&",�H����:�E��@A�'tP�	Ff�}����+��J O���p�[���4/q���	]7�3aq9��"T�g%��d�9�_���q��R@�چ���^t��ϸ��z���K��i"��l��q���%�8B�yYZ�C0��������B�{���Q�O����bp�(�p=�u ?�Xd b!fIf0=H"׾�aW� ����љ�=v]�PW���ʤ��� ����$}�;,��<�ʕ.���*'	�XL	�T�*���|�T2f�T;�����ڂ:f��Av�N#��s��_@[�M�m��<���*8Pox'�U�4}����O^=���Y�{��}́)�}��Q0�vƓ��4�Io9K������<�"Zm�#kV@
�?y���矼�AT<J}˭wjH5�ҙ�-����ᒬ�8��ae�ǣ�B]�ʓ��R��K��Uy|�����"D6�fsW���g��j����%�?C4V��P�&��ԥ�Q:�O}�@G��}%�K�m��b~x3�nl7���MqG��i��H"H;s�"Jͯ	я��F?�O>l.��<^~28�]���"K��y<2�t�к?\t���Gz��mY�ٚ��R����/+�s� ���n���!1�!�̋�}�5��D��}�o�4Xib�f����)��B��*�� b�$�
2<�3�_�Nt�d5u�e�����3���="��sOW-w�%ۅ�g�s�(�mn�tSw���������x�i�J99iD�����-t�~s�95��I��:\pRs��XK:�w�T��2��6lyJ�vt��K/�
���+�/�����/�|Nb�o|�'wO?d���"�C�=W_Ա�jpt�r��[7��Di�����eaP	ٴ�T�V���2�jD�??�i�LU��Ej����?�����t���Q}�We����%��@ �xcw8	����X�\dJ(J�cs�����h~,-�r���r\�~ɍB�'FK`�gK�A������T�h��`��-'X��(���\�
�n!�)��餪�V�QV0x׭����R(}u+��������o�wR�_TD$���FIw-�0����-�«��W�9p�Y����ӉZ�c� hP�����5ml��T�ת��v��p,��z��l��&djJ���]Ĥ�yMMtCCC��'�o9Ҹ#-Y�8�����3��)�k%�lm�B��n���))5� v~�Wݖ;�0Z��OʉE9}^a��䎚*|�Ӟ���z\Cq�N?�X���Ċ��y�+�Ԓ�hP1)���o}�b���h�m�<�z�Ѽ�F"���O��|�q���&:�m��#��o������]*�ݒdz�O>P��魂Vg�μ�w}�~\j��d���:v�s͕ţ��H�A�*c��?Y	HՁo1�sBx�^���c����M�x�������:�"BBA�x�,L�׭���Y�'�����r5�B�Q����8w�_}�r���́_u���z�mN̥�{D�ſȟi��$=e���I@v!��ܮ��dN&ޢ՜�fȪ'����m�\�
�Tl���nu�?�tY%p�g4��0}~����� �R��[*ܦ�\&w��7a�����e�GO�f�c�48��+�>��?0�Ls�*aـ��u�,��+ޛ6�Y�4���d��7p%���¨~�������	�zKr0M�ރ��]K��CRF)�R�
����?��4�O�o�9������o�n��n ��!�9D�+4��4�)��G#�a:�I���	�r�H"��S|=�@z=��h}cv.R�؇r�0�1��I�k������0��M��*�������������)�M��J�er#����bI�&���#�ϋS����K�b+�{Q#_ԫ��\w9|����w�0�V�d�wުW��@�j]0��7������&��oV�xk�4�u����_�I%h�_"Y��0w���~�m��b!�K��1C��+��e`�3���E����|�	��5��EP�B�ʷ�b�`v�������H"�H2�p�p!>�S���~��z[��X�©ߊ7حd�W]Be���u�7�T#�Xs��X#��
i�Vc%��a�\�X�Vթp������?���Tx־�P�?i� 9��9�'�����/�
����ޥa)�G!,ϒmF�P?���$�,]@�y�+�eQ󡽽/0����-�<�l~��g���57�q�s���={hm�}�`}Iz�q��#4"�K�������T��0��u����/ة�}~&�V��N9qs\��oq~��~D�X�.Ǯ���A�kĒ�*������&�V�;�:#�cTr4���܍���ɧp{/����e�УR�Z��h\����7k|0�ü�A�H+k�z���S��ܦjbX�S�KK�����X}\���|.�T?=M����N��o a��@�7�&''Yi�}O=6�Qf#]>�t0V|,��+�y��>�������18!?��Nӵ���d��n���ɮ����2�Gy1��۝�d�t�m��}���s0+���v�/A��}B�mx��JZV��Jr��$i�W�9�u�,��K\��$�L4���bD�Q�,}�Y���E��;��¬l���Ȓ�I����NLFc2���c~g�B��ɿuuu�0�l�{����_L��͆x;~T.��NON��lc	n�*<����\��v��{�G�[��<Wko�����w�`������Eد<l.:��GjO��J����o5q!�m��;~V�;��/�ޤM��G8��#qv�3�<,KE�ȰC&����?Yu|?D�'#R�����Wq#�c!�� ��f��T�a0�W�0�$�)vf9�:ڕQ��6�� p�+���@�&7�5?O���H#Z��WGe��|���؅�lC�n^__ch3��1b�/�.!PEO�\�l�ͷ5��E+o��tf·�"6��P��|��5���3��}�:Z�>uͱ?�|s�:���|���E���)fg�<��W_�z�L���	��'�,�	Z�sף��.�`߻�#"ʈ��!���0�~.m�9�ß!y�c�^m����~Չ�xO�=Q�Z銨���r:瘍�
`4�ߥ�x��1z�����H�xT�l�V��w�k���ZO!akgf�A_է.՛\��'e�B�9^8��b�l:���U����M]�Bm�p��*����^�
e)�o�ȹo&�~
Wj�g�K�h��[�z����aP��Q�@m_��"͜��I�fi��w��	z��t\ ��#q�y��)��+"�x�V|*@�;��~	>�iY%�[%����ͩ�7�NՏ�k�3��hk�;U�5�%�5dv����N�b�737'���`U�wed�m�>��e�m��rs���ZT�'�v��n����Z�%�M���u����c���u��&�z�,�:6�.a��8�nاD�JL-e�uև���/¹+����̷�r��h�غ���C�j	=�Nt��]�ga�ں�v\�Y���.�骎C�GՂ��3q-����G%lI��S�
Y�4�ۧ;�&%�Ƣ\5�I�.���<З\�ڣ� D���ZO��� FD�iN#�"_5͘_�$u���(����0���\T�G�lX�+�p�/Ow�Yņ��s\��"��|�G�/���Y�"x*����j�>|���Ŏ�@�Ȃq��I� �W�o@�������+�~w�� �i�7�%7�A������"�]ވfM��\�>�3�Ưg����ZIz�J{�Rأ��g|�4�UQ!���Vz�2n0�)WT���������P����/�ƃN"�D*I�!���DX�����m%��eX��Z��� ͻ�ܓ%s�%�u��d�u����|��!��aј5�jF���}�E��H�U��^5���i��UY������%%�L����P������'�x��8�� Ɖ��ts���1}�'T�E���Y|���͌\#��I]ގS ����g����E��-�� [u��ۈVl ��}7NN��1|�'���,�}I4L$j�J�����>mM���ʋ�����B'�T�ah����`�$���_���^o4#/�g׀#�~�A"�n�~,1�2r}"`m��fŒ:|�
Zb9�>_85�+S(���#\��0퍝`�pVT��%�w��
��)H�H�w���ZT����Z�Ԣ�]���sV��yGϠ�������"cX�%�SEf<��ۈ�M���ܟ1���|}�]�B��Ƿ��>��}HKf�@�cNW�o����E�������#�ǆe�΄�*�b���^δ�% a费��:
=ܿ Vd�����(��h��H�qY��nYW�� ���L6��P�I���9q@~bs-!xm���*�e�Ͳ���~z�����7%�ۛ���o?�6��=�o5��2�0���O�>�|�� 2�b��1u���W��w�m~����LC�?���Q)+��r��|���\�f v�$����������>��֍9�6�v2#�?�sv�-�l�ڭ����`�7���|Id3I������z�kGߗ��]��7����G���Y��K8�#ސ� �@Q��y�	S#{p�O^>�!$��r��\<�I �U�������Q� ��T��1�r�̀���f��,,*)�	D��۷yVU^������C�
�� ���������ڹ���2}�c�����V��	y�W��k�&��4���j'�x��ဤ�r�m��">�; �-t.h���c�#G����; �*���Wb��ϊ*�c��?��#��G�u,/`>-H�1O:
�(�9��(E4,~e%�h��z���X��B��l���%�#,��+�Jņ�f���8�� ��ԩVV5��
ִ�V��p���_�2�\Q�ٸ��Q�=�򱺥z+ ����f:�)p�����|�eTUa6Lw�$�i�n�C$�Cww
�ҍ�HHw�R���Cá}��y�o����u����{f�k�����e��u��y�(��<��d�X��Np�[�E��T�d	����?��{����dƮR�q��S�\`@4�|m_��ל����=��6�S�'ϰ<S
-��h�<:2-�%�>��Yu��?Q�������qw�i���q��_ՙ�S1�j�e^���%Ӻѷ�D��9M.�P����}��ul��FX�\�����GGO�V��,̟|�HS�ϡ*�Z�2tL�<��'�}���_�����5T$��E����'��[n���i_�o��9�h��<�k�6�3<��6U�%5O<¨[V��s &�<�`/\
�i�b��� `��J�߆�K��$X����y�fo��7ƿ/���n6Zs4�3�6b���Z�Y�+6�Ǵ\�C겋���umC��0Ye
�镯9t���я�tg���k���|:��]]��JA�t�LYbf��n�����W�㓓h^y_�����BqN7�*7�0ާ7V�X���V��T0{:����a���	�D����dm�wc��%�7�U��їgU�	�
��p^�~<%b��7Kx�x��_'���{��U�)�X3M./��x]��ml��W~�՞�[e'<焾��e�dB|�|�����*1 &x<%$�]	)���|ݴ�AZN���t��)����?Z 5�����묢��8��0�DfX�!���kV	��SQN���A<3��"8��5L5�-1�|�b�^Hw�,e��3�l�c �q9'RNx'�
u���X����{Eϰ�J�a�h����.�ϔc��EVJ?uCGiIJܘ2���3Ѷs�ul���M���%����\�=B~U�� ��@V��B�wM� �P|ن�����&hy??�� e,Ff�.�u�<W�ܦ/OR:bY���xqY��3|�o���5��b��d��'��M�rmP�d��>M&@-Ԑ�I�G�|w����~p�YKpӄO,|g5��TA"A��y|y�!L���k�f<�.�͗y���gz�w�����n����.K
�j�n�9�kf�7r�Q$����C�O��φ<�(�3C!f0�헺L�2��R��}ۓ�o>�0˜d��֗H,�� ,��?!PYE5$�3������js�6�ߔ0v��~<��Ҵ/��r������i�1DU��T�Ř�#�zBB�F�o��gRBn������ƽJ�Ӛ>�'9��Fq�'�ѴC�˼���ׅ*�>�!����O�+2&Î'��<�ܤ(>{���r�V��,�q��"�>��Ņ��`[�D��7!���ϓ֬�F��/)�����l?��g�}N��v�K���]eP]��GP�q�~ܶ�I���M�X�c�6�Rŏ�(����Ē�����)q'�Ii��X��ؓh	��D��W���~�F{w���W2?䙂vĻ���z�Z�������V0�!��C��*�u���J����za3��}�����N\��&'�����*|6)��<i�V�2�"�bA�&�?8�� �BW���~lm�+�\6��o2��V���1�<����/�o~繯��|�+��,����R��g���h�	L�\7����8�s�?o7���|��� �+�`��JZ����.�Cm>��/���kI>�n�߳�7�������Dp4�/�^h٠�� .Aclhjv*u�K0N(A?�5��2�u����Ӝ��J�zfJ�vhZ���f�iZ��nyC}z�����^��Pf-�w����1���m��b0j�K��������t���v��{ގe��w�	7��4Ьȼ
߆�OOs����	���n���M5�@�=?3Y�ӭ�&������kc 8<r��*�(:����Bvp��*�
7��혉�4����ަ!oX�is�Q�\�ا���n� t.��Ǟ.����z2�u�V{�Q���X�i����M��=�����,GD����d��PB�f��s'/��v�crjj��l�P{��������w�U����2��NF�1��Y)L_t?�69[ȕ;�`aDQ��:��G�^�����S��U�ݣ�*��P��dY��G>9��}�����>X/O�����͛����Tv� =�7�}o$]廃���W�B��w7��Y��> �|�n ��f�{
���v���������8aݞ������z=��0���b[�\�W}�1��b��L���_�߳k����QҐ��n����sb���X� Ot�^59����#]�T���߮�k'�|.[�uF���]u|����Ng�����Q�̕�},Ƥ��>&�������e�#�>�E�3*�^�-.|����/��6h�������OK�_���K�':�8���p�nڨ����Q�z�(�h)����!g�$+1ƷL�o�5�rot/ ��'[-�S���2Ja��y�<���XW�V���^�x��҇��q$�d� �=j4�|��-��|h=����c�����kjhl;d����CS��g"��D�_�/G�4=���j/�X0�(G^r��]5<l��~I�#�P�ipEiL�����'Q����/
2LM�����%_��C��OG�4����+��B����TM����P����_�p�a��!5�>�N�W�⿖��4@�.�󫈛j����Sm��?N�GQ._~�kyĲ�����p9Sd��N��?�U>]g��	E�(��dJ6$,��ǫ���/�m	#*Ar2����r%^����B���Ɍ>U�>)�Nr��� p�L�N�{��lrɖ*�����2 @
��d�F�qu����'{(���Y{ZW[�rL zr���b��t����:�D�"����t/л ,s`�6�#&�+=
φ��D�'ïuy){��0}��, ��WP��@��?wn9y�?�#8���/4� $M���{�/歎���eH����?�)��7x�޽�o���g�	O���z���+��S���䁐q
D݇wE�0x��NBp�!E�Y�O�c�N}:�E1�g�$��m�1͸5�
ޤ�Y���7.��Wl��&����W���D����������z�5	�c�m��1g�c}zi~>�~��t���ѕ/��{���Vo�D�K+����',z}�v?o��,bwdќ�N�Y=x4ǮI�le�4�5�~�����C��֏���11����;�s~����"��|n��J�� ed%�Sâ$/yO9n=y~ZF�X\I�齗k+�4-2!W$�´�A�V�G*~5�,cY��ݙ���{�*ġX�~�+�����G��3D\�P3�����/�$_'��#"8��q��� �i��ܰ� �1</@�VMc��~T��g��jy����'���g;Pa���Y��%�Z >30<��i5�����!kK���MUt�<�
�]������9�h��}
נW�8��qҖＫr�:�#5�Xb����pV�U?5i�ʔ,��e��c�y?�����}�ȉz�רZ�'�2ؒ��?S�
�BZ��w��q�߮�-U�(F�+aӶ�E��5&�����|��l~�M�Ǫ�vz�<ն���&��3>��
"��������D��p�a,v����iA|999p=_�/�B�,��- Ɏz����k����O\�ݧ��(����&�t�C5�A��%9fb\ae�d�������-�R���r���ѥ<:O�V�u��N�z"��}�	�*��bλQ:�.�����`ko����u> �s��u[�[�׏l��wg�MM�x��O{���YV���ވ��SfYw�P.�
�v�w�)њ-�ּ�z� �X9f"�:� Gc6��N�T��Z�-S��b_֠Aj;v��h�?�bH�B)D�`f�u�p���M���PT�D:DM1�7>(�z@��kX9�76�wjD?o������ԧkP�HxJZ�zݫ�%|w��g(S��O������x�}
4��#,|��@�`F��h�YW6"����Q:_�ji�!�ó54��l��;[�e5�j]<...��#S<<<�}�"9b�.f�]�#D�������1����(�O���OY������ƯS��7麸�u�6��#������S��)���F���Q�Ϟ��U����&�L;�̼u�/:^㼱y���jX7 ��,�X}�m�}����$�;��jm�X�s�8�����ln��'nSv^V@����vӧ��l��;Z�B+%���R��z���rX��C�����7��%���,��x�>Z�Y����A�bWۗ���2j]������k��rzw'�޸������x�\=�d˧F�3�s[t�tg�q���9n�,q����D��:�����M�l�_W�#�:��<��ӴD霹P��`2�u||iyYE�n�sI��Q2����H�+���:�nc{P��~RB0�w�<2=;?��?�U@'��s�m ��'ͦ���XQB �MTj�y���<;�s=��k���Ч��sP���v��%/���)�.ki��-��>��r��WZx��
Q0N�����=��J���zF��hԞ�|��ۭ����^@�6����O��a.��Ŭ��c1���{0;u�e�,���5����$���	��䋋�T;��n�]&-�*	�L�����ځ-�j\Ѫu�*�� @^��_�:��P�����I�xv�>Z���Ug2�l�f����/��Vu2�[8)�ql5����8XX��s?֤Bcj9կ�6s߆e��|�_��;������[�BH�Ȅ���!���e;�~��O&ޚ�;Y��c�����/?��퀯���{���Ѹ"����t@@�¿l�~ߙ�����i�P�ceXJ��$>K� �,~v�T������\�Nt5�m,�0��f���q"z,��X�K��J�y@���`��!�J����Aw���6��tt��,�j�Ƈ�ŋ�r�[i���zE�EnRw��P�D��=�����!_I�d"��T���""�<#��WBN��=Q�eN��X���YX̴7�}�@�*li��FQ�#��7Z�o���#��W�-�u,�S����D
�<�g�no��`�.�2�5���{R�T�V�~��9 �Pf��3B�L�}zz��qjq��p�>auJ�=����w8^�6�!�+8o���K��(Q��ag}R��hk���c�`Ϟ`�^�� ��Q>$0�*�>���:1AQ�W�q}}�x2�/>6��������8yT��୭���,<||��Ck2zUY�[��<U,F�q	�導��Ƴ��lܰ�.���RX��Y��<��`y*�RV���%��}"�D�׺�|��R�b���qcXl�-���k�w�bqryMMT@�;�,4�9QX��D��/��}��t�@m���˼O��s���&TP.oL)�a�C�;��h,�~�6�Fu
���&�.�/�O)�����؍��$�D_��cK�`���4S+0��y��Uf��Q���h�l���$�҅rĽ��uR�w���|B���lu�;�^.{@�p;�:E�?���i��V�ߌx�U�1������I��1�j�!�)�]�3���YP���#I�j��eNV��7�#�h��Ԏ�|���5��h�t����$�(a�u��Ky����`_SK�ʊMTL��r������p��r��lи,�_����F����YX|��87UU��Xk�gՌ����Ja�f��|���סMKy�������aT<�V�T�L�̞2ΏB�?���[���{�%�w��S`"*7��Y<��J� ��ayy����6y��/�)�ttt������:M�A/H}��G�T�����aU�x�*!C��X����
~-��pՄ�V�20d+�@O�Q\�M���C=�A��D�&�H(�&r Q�˽C�|��NH��7Yx�I�F�D��k�v��ז4���IDŭP}ʲ7x���`w7;��K��S��H"��|x#���N����$p[�o������b]�"N[Q?���Ґa�z����"���Taʜ!H.�[~�6Z��P�c�>5��m��E�Vu�5r�8����C���9o�����t�p���,���Z�>|�Lk���T+N������ؾ{SW � W�Sq��7�`[���6��r����N#n�ԱAඬ�`��.V��ÚĮ��>��g ڃ2~��f�U��lB�iM~�(<~`�#���<Ԡ��+A�C�
�2~�st���f,r�a�=gDi||m�f�;(Ң;F�f�=�~�K�9|5ۼ�Fb��Q�(������3K*�X��&���[�%˟g���U��#�-Ǜ���.w�R[�W�H座&��===��n����Z���Q���;t|��Xi�9��/�䲍�h���~���w���>%e�:8�ޤ��"a���S�
�u��5���WGK{gUXD��%��/�=z�M	i9Vҙ���P	ƻ�\A�搰n�k�>3k�rhXߤ���������;�V�*	F�����<���iI�䪢"�Uf�[OmV�1��k+%��Ye8��ȅ,������g�T�Uϝ��\�ŕ���f�:-(�s��(y�jN|������O�UΛ�b�4E�RE��em���0�VnK��ػ�s��=��S�ӛp'A���Qt�㭨��jِĘ�����;��_F�j,���C��{���;����N��^���^��
|�w��x���V0b��A=Ekձ%c�L�b��`�%318�����@m����i�B�%{�ZZ'ڠ�����̟��6o�����UNN�%s�J�[Z2��.-UӚǡx�P,�.�}��_��S��wA�pX6N䠡 ��$�V�;����q#f�%��n}C����.��ض��u���g���w��bi�jo3 �c����I��("�/@��s������6�^ŭ��8�"/eo�g6>Aa�7 ��ir ۃJ@� �d��_2J^_��]\h��v5���9}�	�{+D8y0��v��+k��YO�8@׾�ӾJ4	�u�&�I1~{����-��s ��y�U��C��\��@�T�J����3Ȏ����^��yE���L ��lP;�8���{�i��18��Ih��\�_y����DC��`c�7��<�����[��@G�򖊜2= vZ�N{�4���E#>�O�#�va	�ܜ��]�Ki�=+c�/����w���ވ��G�'�7[��
�{C���t�/��E\@>Ń&{yw/��j|�W�xL���ϴ�e���ǨY�P[;����Q�Lu8��A�C��/�Z�E��y.�,]��ea����Y�2n���Z��хU��/�Cn+���'��8e��m�A��3�F����IB����y�6�x3`� �;8SHw#���Y��Ǌ��� ��ʢ��<b$�At��2�K�!� ��D��OȥNt aNP?_~��qj;���d���Ťn�V�ex�A�Ņm��S�����j�s[��橚�� � ��n��=Vs�ws��Ǚ���$Z�K\^�[w����R�K5w����˼;a�vc�3zS�8�룺r�wZ]Q�A	�	���Os�L����U�q5�3i�h5��Ldx����G�ֺN.5���+�����ݠ  Z�Ƕ�ܷ@��SaS��ٸ���O_5��x�@�(s̻z������43�Z9J���+y�u�rBڻv>�/8�VDx�Iz僜�i0�r4��l_�c��0���WTV6�u}�H�R̪�wĿ���9<�����W����,�`$��'RI���1}p[h�UǙD�lg52U�JdMud98�t�	}�DQť�����ag�6Y'�+���P��d=��\��&����w�jp�=8��ź*?`���:v������t~go3=������=#��4>�mI-g��ӓ������>"·Ԇb�X>]��z�O[ ��!�M�f�"�����'��KX�I��u%U�'?=������V�t����d�
��ހ�a�~�����(���\`��l����IC
m./��ס��3>>��}�~����x�?5�.��S��8߉��8D�J�]�[��0"����/j�P�֟�돊����W���Z�TXi��Hs�w´�N�_����;u	�	��LLL�������
a�AT�/??�*���B��
�w������_D)2[��]Bf��>h3�ե�r�Ԣ�E����V���um�Qψ�vS��U]��i�KC�y&�5�� qͫ��" '�q{��@��o?+�Y	����8����#�'٦�ǲ�4�ػ����^/����.����3l|1��@�!�~����n޲�� R$�f���?c�}R��5�;�Yis�8e�݄M--� X�ˠ����6�>6��5�P�?r���S�<����d��p���N��H�U�Wc+[{b�2��߯�(M�^�Ri:��3KL��R^4�H͒���(�~�9B�aI(p�����wz�!w����4������ [!s��m�_$5M��Ѭ � }��QIĞ(|����g� ��|�p3yp��w������Ҭ�,#�E�dZo3A�ë'��e�֭�������lX姹d*�b�/�ܧ%ˁ=z�����;"I,b���*�����P�{�!��8��b���@���ǲ��w-��6%']�b�(#b�=�V���C0�����w�o6~kѭl��O���k����v��WVj����bU��Ѓ���q&� M�Ծq,,e���.�'��$+��6��CT\�¤�V��l�
m����Րq~[��6%�X~�I���d�/�hx�"�Z�t��{�y�2I����@Mw��J6A��'�����j��Z��p�)��)"��KF�[���;R$���X���ς��*U �&2���8�{��C�ZZ2RY��/߼���9=}lf2�)�r��tn���=G?�^�G������א�8K�2}�Zf��ld���X����"�2������S��wD��ˇ���T��k8�3�����cV�(����y{<p��s8Kj'E�p�e��G���7ԒW�TQ������<!b;���Ō�˩w8J���xv�g�Ծ}���?_L��;��Z��8I�;�bxz�ȥ���I	��	�(���k�)>^X
��6?������蜌jS�Z@��U��@3�!iN8$*��o��-+��\{�p�c�V���y��ț�6c�w�qO�^M��%���r� 1D�J��&3���^��i%<�:~,���"�.M�>�A䲬�|
�>~ȏh���7и3��jҼ�Q��|ںrm�!X�Tӹ�[qY���!�߽�� ��n!m�� ��ht>�'%�F�L������	�����:F������WxŪ*�N�+��D�e��VNn��WD?��M��ʪ��J,�W8v�=��ܓ�2��u��]��>`���6"F�&��l�=�xd�A3.���˚Q\$xd�
F��8x�__���}%L���H����Y�2�f�tq��J��GO(�/��L�$/'��ʞ��z{��v���z2=��wY0��)m�)�P�X����D
��.��?+�b$��~��������p���������K�ȭ��b��#�kh��[w3Z~��-i�-��V��{G&�4C�۱J���j{�*�NE��j_��2�t�V�XT����_���|n4��۞ڼ���Ӆ�w���@
T%e�@8��]��*(�Z��e�yYM��)`��I�r�8����Z��JX%�9���DGl�y짬��[������ʹ}���H-�m����ɷis��{܋�}�U%���}d@e�9��۱��XZ1��2�;���0�og�ķ2E"F��Ix}-�T����F���޳`3�B�֓WM�(�~������m�5}'����_�߱wO0qʓa5�	�nps��枞ׯ^�yq	{�X�|~	�U���J�h��V�f[���sa���w��y����]/���Oe���P3^(n�Ɍ��/�6�`�u����&X��g���)	���`�'�!����v��IMg�$����	�5����O-l�R��U��1��f>�Q�w������V��f���`)���`�&�����v�#�q
����Y1��,z}W�I�.�m�Ky���?l���*2 V�֣Lx#s���@��~5�v�W)DFG�GH��H�_y��L��ޟ�kq�=��p��[[Г��>Z	>�;<`��d��"e��|V,�y�B!Xې!�Q���>l�}ơ����,�l�uܟW��2��� �"��E&ZSb�/�o��V�9}%�Q���S�����Lq�����t�@��1/L�:D,� eߵ��|���YZ��f���|�_��9�����;7���zn�~5jN�0_'�b
5K����i����T{�0b�o��v��@�*TB�,�1��2:��=��hɯ_�x��5��(I��zg	�?�ZS��l�4�j��Z�ɗ��[����d�1�8)f���7��?�R�r>��=ف��3)���������\��W��`���Ad������w��/��w]�/:���għݼu�B{��w6c��Hr���>�*����}��$s�ٗ"��{ϣ�4��@��lFF(�k�Y�D��u�s�\v��fZBl�Sm�wpA=Ϸ���l�g�hOо!��Q������)�����I���*H�������D�i��]�!�хO心��F��p
i�� a�D�W,B����P����2��Q���R��Q�~d~{�e�R�Я�'�ML1���-��z����؝4E�D���(T@J�<v��<f��#��{�kr�mK�e���&��%�4�w�%�"���	�F��M"r�T�gxʸ�?|ѣ�3���Z9���a��.�b�U\��������~J.� 9*g�y��q6��K����U��2��&�G���9biho�����?%���!^Aˇ����^����lu�4�YO`�����O��
x��������ۮ�:󛗟�2�ajR9�ͳ���%�
��SL�������Ir��k"Yc��\���`6~����κ�U	�,4�ʆ�c���s����d_���M��|�����X��/�J���բD�y�7���۸ﴩ���أ�Lux��������x�2��l�j{^������(<��R�@M{�a�QR�/z����l~�|�6�����>D�	Nb@JO��r�ui����S��Ə�P������<�&��oL0���I0}���>{�U���K��31�_@�3ʓ�v��-I�%�#6+���&�U��j���a��/��\�*���J����m��\t��T&��㏱pL�vrc;�Y;���#�c�2Sm���o ض�K�����a���"v`=�=p�7���� 8+~~�z=��V�А�a63P�yM�sq(��ny�Z�����=;i��[�?�����Q���h3����q���Y���y��$l�֔��_��L�.�D��M� 15�ڽ���bd�ǿI(�^�#�����\u�e]9xr�0j�3��LG�Qb^�
ݤ�dt�ʞ=(������&O@�==�߳�`e��?u�mߛ��~�iCL�}A݆!��҂�Q��	*$êߵ_LX��4��6r���Ծj�����H��o
�խ��6! �*#� �N�5%WM ��	�
���_w�/ہ���f.'G��|ZBhj���������P��x����{�ygۤY��{�G��he��Pr�^�	AKK�q/�*x��I��^++㶟f���H�;�Z��f笭���_���Q6�����3D�'�8�KR��X�4ʛy�CNi�wEE	�(�x��>ʅW�����t� ]q�]�JR�ۺ�"��qk���-���f�<�dg�j���?����4˗�R�n�?UA}{W�p����(��o�����?��F|+`DRs~�o�X���;=��k��+�?M|a�DGVf$^�\�`�=��0,�%l wQ��b���Qr��-[h,�!�����������-I9@~�­<'��\��xț��ar������"��G`[�W~)GzFF�� �/��qO�^L���_bk��&�
�������H�Fx_��]�i��9	��}ۯ9�c�c�pK��@={�8��K����~��v��qƼ�ֺ�Ož���-|Q�a��~qʭ�6������df~�A��^��mR�rQOՙs���'��x�<�!�f��ID��<]ӯ����tB��nq��Ч88��i���S��$ �2SR(Q�6s�p��u� ���Đ���S����yp;hI��ܩ!��X�U\p�ξb��og����c��l����1�J�8���W�Y�@�Λ������/ځ�Y�b���VdBz��h�,�HX
�B�/����QY��+�=��t�K��tUܟ��&^i�ݣ�j�.{�T��b7�	�}����O���N-,v�z^��u���u6���:z�ôs�����A&�ǆw�%�YIqV��=.0���(�� g��|�����a��foCO
=X2C�5ɚ�2�YP����(�Vh�/��$���!�!G+�1@(C���9oX�n��:ID)Iæ���X�D=�m|\�����s0�2|Z�� w���J�p�a����� �(:..._�k���̓�j�]e���W��Nt�t�p�P��?�����Bi�S^�0�Fr�d�y<p���a���Zn�X�*,J�����ʕ�T��?�O���y��1��+Iw�j�ņ���?��>�եd����WUou|�ۓ?��p����)�!�l��1N��o�\��)1�m�M=�±���ò�4�����Gp�\�@a
�i-��|���PxӨ�c˴x�O���-�-�7�^=5%~.���	/�QW�M}���	i	�����ZD�缆
-e%�C�m2C�ƺ���6]
�<_�J��ň��oU��@�b ����ye�G#/����mP���E:bø��L��S�x�1�e��is2A�s�U���C�@	j�vɺ�xu ��1T�E�E�5�����$����$(5A�؅����������������p5M����,ȏ۪^8��h:q�:Y��&� ����b*�{��Sw��xCju�xC� 8�N�=����SO��������1p�S���,��G��6~J��V�k>m���&9���ZTbF�2�2�V%miQ䖼����Z	}�x4i-�����I���8W�3�&���U��z$Qh�7�����TY��n�Q�"��<��Yl�A��G��M�l��_m
o~� ��&������<�4�����	U[]�G�_$g|E\���EܚF����*6c#%�)o~��f��a���l�7Aԋ҆������r������̗�@�=�Ç>qj�+I���M1YK���W#ÉG��
��m�&k,�9n�9����5��v��X��"R^hԷ�v|y)���:�>+�R����A��=��������y���z���J�y.�����0Q~$�s�����>L�F/`�!���l�E2���ѺJ�JEӌ�Cǩe�����D��$8:�����͘]Kz0~�)��Ŭ��?�����u=��CW2�ه��G7���Gϰ6�/�o>��]��j��%��j5��F�M����]�.��$�u֠��c�����K����j�7�2#'٢���LIK?��g���.��@�ՒZ���c�5�G�HV�J't��ilF4i��� �5�����S^B'�D��/Bìv����'� ,���m&��m�C7�9mgy�X �S�Qh�p|���v���쬫G-���X5Ҝ�5G���$��2���D�l����}���)$�Ȳ�Y�\;�(�p:��(�I�zx�;d���<N>ȋ�j\}�_<}�z����kQl�8e{eu���!��5�$�׻E�9A�D�����j�^λ$��O-�t�܅<x��˜y�~���R��[\c#��abܧ���+42���J��/$��f��<P4�e���\�8ON?j��S�3*����5׳���z�˲�kNpCQCC�Wlu�@�/Er�U�p�l�lAf��SEd�o��f�q}<����H&ِ�Y�6��~i����mg����	-:_w})I���dH1i|].>'��h�L~<�x�J��� ��UBv�.���z�1J��q��]t4N��q����v��'�q�ol<�Ȕ�@�v����^s�<Ӫ�KM��-��2@t���[8/n���H`鄑8j%�З����(��]��P̖d��ِ$1��U3[M�"���<�R�"Dr��}��I�u��]:���\1��%���1���sP�Z���� -ʘ�Hw_̼�tZ��|�Wj57� ������ ��M5%�BP��s�M+��&΀�)����V�S���=��a�R�{`i)�ŝ��-:^O'�u��?�[WGfhh�4(�ؘ�4�ǣ1��{�e��W�Ѵ�&c�Ke�i�D��'���Wa?��_�(`9IczȾ�V��1)�L\�B!���*snQ��>h��a�]cJRkE�Pي�D?�˦�ٙ�VQ��>=L��7�W[���9���!6Wz���'�Z�wM(�j�7s�MٕRY0��6|:9p�Y|��O%?n���Jg���i>��<���zB/Y��J%�,�缁;r�9�y%[=;��~���῍:��5���I�|����A@��p�����AnP�<�R5(���͓�G��.\S�y�H�f@�����L9I��8;94�$��ˁ�Vz|y��r������v�	��=�L?�cυ� �Fi˨���^x34j^@�o��!�G�j�	E��Ȣ,��*VV�N��z���q9'�(DL*��v'X�CJ�T��G��SW���Ō���U���+6Y����[7K��>���k�iT� S��t{9\�����^�r��r�0"Q�!����ͧ�$l.��3�E��k���	/t�2��"���a���d�`z����mL��(�{gW��~�l$����>Zխs�U,���(�5MQ��g��wy�q�E)������F��Mt��U��|����I\پE
�	L����N�zB�{��n������C�c�M.;����/S;;<p��1)|6<��%:py48F961�FL�~]8j3��փqW˪`�|NTggKv�T�2^=�8=����������Z���i%$�c���G��v=�zihq	;�k� hs��ݚWE�S��5����\?>v�q�҆�����J�*��(�"��������C��3u���|���!�/)�5�q	��[��VJwf�s1�1�,��d~��Y
پI`��2�_M�Z7���!7m��V;��%�F�m/�G�0{����L[��@���{��;ѕ�3��̵+7����vA'8��'ײ��>����4�� }V�RC"gjH%~��[c!�nX�xρ���q��B�3�n����̺�ϐ
��;�n�i�1�E\�����I�ͧ֑��@l��^��	����L�I��88�[V��l�r�]�BZ�.�*C�h��gK�6Yn��,:���O��=���l��\<F5�)�=�g� s�����3:8}6O=���N��?&՗�����*,Ϳ�lӪ&��I�Ƽ!��|ꑒ�W���I�*J94OS���.d�R�5m��{Lo�;�h��X�,#)M*i�i��F�頛A�F������Xl},ON��l⭁��Ėo�z�a,0�1��/m\�����<]��6i���.���}��d��.F�&팸:�\���*	J<�-��7��D}�R���$)�A6�FM���u%����Ew��.��+��eO�:�&�V�OjQ���=O~���9n�Y1A�x�R��/2�l���ُJ�Fڝ���$Ɲ�;��;�g���A!���q.
E=�A\Ҕ��(�mp������٘�m嚻���4�_ȥf�/F�jx+�����\�졿�nа�����6���C�#�<���v�ZX��ɯ���U���l����D#�g����i`I[f^ףl�=%�Ɍ2a�_k%�ӫc��ݬ�mY܅'=����߼T)ר�0���9�yg�����%/9����%d��*���7�no��/jrVA}4������V�e;lHu�����1L%z���$��E%ߝ,5�bU��[�T ����c�~%���-c�c=Q"��8):��ğ?u3��AA�f���⦿Y��9��Z�Nt��5�|��8/��
CJJJ�'�7$Ǯ��E?��ywV0�e1I;+�I	��V�^����{�5<���Qy���a�=�Fd/��o��Vv���|�1��xo𔺯P��Q���L����y+D]^��-��^��S���V��k�:̅��ւ���l�`{k�h"�T��@> @�UP�XW����G{:���#�3WG�Y���{p8O��K��?�+�W�R5̻��;�X��-�X��_���Z�i*���ݝ����jqn%���	('.��M��2���FC��FÐ�u.���rt9��ye"W�:p�
�UP��~w��Ck����VB
_Ϧ߅�
?�B�m�eQ�0R4���r�,_���@2��S����}G5\לM�1>F����6����X��6ʁ��V�w'�M���z_�n���i7������n���Sb�����n�Ut�jX��1F;���b�����|��n��]�s���&�)U��piƬ�����YB����k~�����<υ"�L�����ԇc:�}#-�d6ߴ����fv�h���ܹ�Ff�P�HǑy�v=��S���h[��3uR*-�����i�J��5r�J�}D'�	���d/u/�j����(��v���3dد�ã��˓�[�*u'^���2,���A@J����	����$��n��e���A������������.x�㬵�>k��z~��yI	��C�iD�RY$�bu��ܜ/"�/����Z��e�o�қ�lM>l^i�,�ޫI>�ն�+�ǭ�����������6�j��o<=?����\���dp^��쑖Ο��]]�0���T�z"D���|pP�����5�^��{w㔜�6�@��8_T��
�����=<��p�f/����u��;�U�Cv�l��\3:cxؘ&�B�;��͑��������na9ws�qG���J��bٛ�e��n�0/�(�dqG��H�`iǐK�n�����p��Y�I�L�XV�2�}�0x�Nm<�.rx�O;G��;�j�!"!�k+�~݂�0��xU"Y�E3�kx��81���ȃɹ,"
m톶B�1���C��s]�j�|,dh([��<�:�7QV�CQ�k��+g�$O'�.*jy�]�1�t�1	�_x��߇p��y5�[�Հ{G��z���|7�oC���!�4����C�H,�a�kļ�V��3[*��J��~��3a&�����7s3��
w���җf[�!��YL��kD����ܛW����i)�!0�r��is\pMNE���gjP�ýV�7�}�U�|�]��j��&�m�˰`��u�X�ڱ�G>Rz+�Fc'8ϊ�:s+ۛ<�8p�9A��ڛ(���Af��畾CeY�zw� 0F^�4|�N�{�y�T*qlr�%{�V�q)�:�(=����yzg�F�G��kJ�P��K�>�v�4Xd��e`}6X�Ou�7��g���7�VĄ�����&=�7�����K����<!�'5�a��¤���o ,]�����C���3s#���7�{i*���� b���[b���o���hW��PZ��_G\#&�̺��_�/���mh�6�k�}�	�7g���`x!Т2�Hj��!��൤��m��+^O ��E��$�y@@@���F��y�ݟ�rQ>�hiko��Nԉ"��<�����R������0[�;0t:�����ygR�,��W)J�rka�?�lq���+��������T��"9����o���xB��j�sG����ׇWs��U�4���HJ&��E���:�E����w3�#�c�YK-d9j1�S|��[g�J�w�֏�t��!S&�.H{5�'(�"�r=��D���!��4po���͇�=�]�q��13�aA\��.�;�����>�'�e�k뙧�� ��uE['���7
B�X�"Ja�3�1b�pfWB�p��p����Aw��rS�k"�˽�$��r��;^�Bu�2��h��f�D��ui��~��C�B�YI�i��@
# /Evx��Z߰WlӪ��=X&|���d |4���9�$U���W�Zi�����I��y|� ����pv��,�0h8�n�.��n<d)ȿ�����yJ@J�)Db��lw����o{˪tX�8\|��C������4A\c�����Dm%H�Û��%�y�*�<ǌ�<*`�K&�~��y���L���Q���j�����|*iG�<��H��E"%8�����C���	�	��G[y�V��C�����,P����4�O#~C^�(�7��h�q���Z���a�I�)�(������c����ɼ�ɨ��-�W��pW����ڊ�_g��2r���|�� �*[�����7f�c��Y2��e����If�c���T�-�;
ƛf{2���/��2�-���yuY<,�Y՘�1B�3,��y+`�	�e������;/�xx�N3ws���h��B�,i��c�\�;;�&! ᇱ{�GS����[�j|u�Gǚk�};�ܦ�<O�
�F���=vRh�)��M��ᱚX�kҟc��PжR�CKn�2θ/�Q@#}n��23�[�G���A��68��b��L_����Ӫ��d-5�A�2�	�Tϵ߿��ՖK>V~LđQJ����<9�*{�^��|_]UQQ�%�� �0���Y��'{)������Op:�����<�����ú��y±��)�W;��Î_#Tn�:Z��t�
Uh�I��"+������j��$LZ���\j��� ����	��?Ə�9�kMn_�P�+k�^<�r,M�]�_@PoB��qR�DA�b<�`*Lb&|?00�<H�^?H����k���h�:\9�k�e�����z����p���M�Q�����v�ͥ����Oz�K�ٺ��m�׆o� c�$�AdS'��qӰ�&��X:,�o�A�IfM�F�-������%�,�S�!�`����0T�T�Y��D(���'�!��S��ي�)y+�gA��ݖ����hH!�ċ����Ra��h����$P�?C~���Z	DX)w" %��N�*��H<3n�A��11nƑ��k9��[P0��$Μ����#I�]vHcӳ��a�����X���E���<����9 K�U��I���r!ޔH��n�4�+S@��7^?�q� �6L����3��p��ǌ�q��aG���F=a�r߲��2]ei�ql�1s�	����v�>��"���s#� � �,�YYs���������dU"�Wo[���WRq�L%$n�6��xt2��$%#no�`N�yq�!<�Z&z�6A,���jc���
�%��+crAf��V'�͢^j<�e=��_���P�Ǵ�B:���d���?��o"1�/q��q��ҹb��kJ���{$V��ͫ(z����'O�J�M�[��*'4Ī�� ��� Q�BlT�i�5���Ս4C���+��a�>�k�"���S�P��ZւQ�j���Q��y{"�����w	�B���n������SOS�(SJXE?��iy3r3���3�a8���?NQ(�ԝ(�YW���������"x㹡�Y��G;[�F�y�~$Q�4�5[<��^����'�������ٽ��S���x�S�����K}���X�����܁�N�;\��:��a�#����<-M��,�E�^���^��Z0T�����= ��ZZ�����֘rYE�cȨ����&������@4����������;� �p]���oL�6�8�q4�414"��\y�<6k��yjzm���Jy�~6��C[��B��~�8����ʸ���{�:o$�1~��k���®�D2�����!jV)��Z;�KNX��Vȼ��x+��V�)���� ���,� >���뵄�����(!�� |��u���%��?����^��¸�6��P �ڋ)4Ԭ������)zªG>JL�SR{\{V�2+�~,)9�65��{��W �lEUU��"Τ�椮wt���H���Ep�cZ����z���f�o�+�O�9�\+�ΎEI}�>O�'�e*�ij��Q�P��Km�� KZf'5�ہ�'���π�/z]-�4R`	m��뛟e�b>�'��a��|$�u{�X/m��,A>�z>���f�<ޟ|���{;tN� 	����Jf�ۤ��UV�,�窫���<� �NkV��I �5�E��,Ņ����x*YR�2`vG�����me��k���0��~ٛ����-�S�f7K:5o��[�:��>8���p#K��\���~k�L��\w�1��
�����4��$�|q��D�S��2���m�o�TaNE%k��]�eҀc+�o/*�]#sSѣ��tF�WO��<�&��b�>�av}���<��R��E�T����q4b�;<P�ԉY���97K]p�e�o�_s-T�c	�}��%��b��8����,j����z\�?<�?�����y ���sv�"�b���;�8���;5Z���a�w*�f0���"#/��8
�A�'�
	�{���4
�������-:��I���d�(��M�]�ɦ]h�Q��-S8~u�(���ʓ��Y[����Z�L�"o���I��w���ʾ.`ބ_c�>Q���L6��!�c�B��+��3Ǳe�d��w�4��Z�Z?'�3[�Ωab�j�zQ˄��d����>�gK�43ߥ�~n����d��OLrk�(��ȫ��I��ׇ�?�"������y��x	�;��۵tXt���f���$<�D$|��s(�f����v�roez���)z���Sv^�败�ʗpv��=���+�%��ǭ�h�KLu��c������� Gw���YB��|*
��N�ҍ������q˻�S�M��n�dٜ;0�P���;�:o��9��<��*�Zy�:<��?�1����H�Y����mM'w�����2R�D{�u#����\������B��n�w)�zY�/bu�3_�Uy79'�{ﶪ���Rc���������[Φ8rb�$���'W�~����P��q.*R�����c�ڳ�G����Z��2h#Y�����=��T+�Õ(=a��kzrA#	\�@!�z�[|�^�60��~��a�f�"hL��R��o�����>VTT(f�	�J�m�B��yr�/�\w���i���G c��nC׈���ν�M���B{��X��ޯM}j\2S����ٿ��_�kcd�:��g��ml���S����T���qS*G�v*Q�j���]�q��uY�;u A? �O6kDA�j��ﾉ�d���q�A7�<�ڜ�Ja�����V�i�Y�Z�:�]��+�S:��Ӊ5U��S�B��q[l�Ta~���B�S��_�n����|��5cK����j ���f/  �5���3ı��;W��ؘF攽��_������YX�d��"�˸.g^��n����ŋ�{����{F����xi|�Ъ��m79ظbXo��V#W�����1^�=x�ΰ�N���O?uu�C �2&-��1�i�c�c��Ăoo7����!UUU�Qr~-�_)9����s|�"zᣅ�
f~g1&r\D��_��ߥ�w���GC�'02�iǽ�^��K�ra��Ҏ7+q"W}�m*�@D_DF`_�S �si�J��R%���Ɖ}�,��e��u�n^�G/�åN��d7Oם	r4�tq�}�j�M��­�0��-�I�����7lQ5�u���D��lGD��2�p_�0r�Kԯ�+��f�Q�e9�v�-œ	m�6��B�����/��q����ty�\d�Qo���D�r���s�$��ڔ��@���6	~������Oh�Wh4�(��0С��}'31L�깋�����[3�,ֽ׷�O��Sb��
�m-��B���O�||����g�2tL0b&j������f:ݲ�۲�o������o�"G?
ƅ_T� �_^!�P�h���S���>������ήO�Ϩܡ!.\�2|�+��(�����46�k�⦻���l�vG�VF��0ț��gu1�^��0%BR��W<ؿ6�ݢ!��OM��L���J�)΀�.V���������A�'�� 9� ʇu��!��\Z�Z�'N�.�$p�遧��Mmq��}��U��"��i�֜_2�6�ܓ�x�,���C��?���U���������V��Y�2�K<��NM ?���.\g���7��R�Q��v��h��呭���Z$ֿ����un��[W���@��T�q�|���-��=k)�C*�|���")�G��Y���9�3n��z�$x���D�o�\�]e��fQ\L�g.�}���(�������k6A��R�ǝ� ��ϭ�$���hVu�&��V�#�	��A=yh��`�C�/а�����o&��-�!��b2�Ȱd�x�.!hJ���o�ı~���nL�hg����sQ���O�k)�j���>\�b�lki
+K�٫~L/��2T���=��Ǘ2����ug�Х��6-q�� go^��A��@/����q�9�2_���f�Ӳ�� �ji��u��v3�=���J���Np�����-c6�K3�_t����R��-�c�����7FU���Eh��K:��G4זS,F����DE:�a�3a�#74��}�b&qR�N82�š ����?D�wR�&g��-;;C���p�e�h�2vgg�V�"l�>Ss���s�S�r�y�K� ��:B�����R�ps�Z������!��_ݽQmQ*����u�����Qoc�J�e"�(k�d%���r�����Z[[3x�������r4쮞��D��S���I<[�e�d�1���������SD1l�LΌ}�
�|c�d��˗��Zz����	?�r�<׸�/o^��c�r�F���f@`�Bg�$*�[>#e{�,��"��U��Q�#�5��"�5Z@˓ �`�k㘽%�NБą�cS��N��[��4��|����>X\{7�D;%��8W4?������/���B@�psC�A}��7�������"�N����_I"x�yP�>��!1�������ڻ}JN�؟�ڐo:S#�u<�ӈ�h�ϵvv;�L}�Bծ�66B���k�4P$~�E+zM����9�2�f���pX�CW���V���q�����gX�����NEnw����90^��1�2P-�x����Q�8H��ژ):������bǉ��;sw�^"a��ʨ�Xm���-ʳ~� �GB���.���d/�)|��I��w�}h�gr�g�KF��;��=��t�v��ţ4�W����DI�B��,jN��B��Y��Lmv���kd�=�W��T<C"���/���@�# -�y8���1su���t7R�8�+�����{W������,�,��H'�:ﷻ��w.\��m%�a�T����g��n��1{�f�{I��v�7�^���}^�z|*& �t$����hko�;����bἎ�����Z^�c�,������f�'��� �*�7,�d��)�!��$�@b�j�hp��L{�#Xkldw3���$�..^W�C��L��e�S4�h���	�����{�>4�gS|�SN�M�{W�ۯ�[z,�[��8M�a���>���2�si��F��.v���T�5����$V�k��a�G�=[���͍��B���V����V!G�W�؛��e�a|�!�X6!l�����}�"���!�hgWU�M��L�-:��F���>�0���t�2��~ReEA��|��C�w������:��!+�qރ]6Q���Jn-:�2:�1��xa����5xm�R�R���_�/ϕ����St��W.��G���֭r�_�quD��u���`)/�A�����ۘa)�I���������i<��q���
��e>i��rvs]�P񥺷L���(�:����3��B.�������T��ܒ�	������0�����`�~�˼�S4dG�5�!��f�b�{��ƈi�r�?B�ܳ��6_����4�{r��;,.r�sw�I�K=OѦCb��E$(�&�GT�Æ+n!�dF%'�ߋ6�L�<���gӬ�ޟPUR����򰯷^�G��I��1�<���a�X��>$g����rww�o'����SV��½nlM�~I��_�5*&��9m'�{��C��|~#I4V�'P|�J�G�'Bū*�&'��͞�ݱ�,����%��G--�Uv��PL�~B���a%�&�� �,A �h�EԷ���h_g�MKT�ط�:������`)����Q��l�b�k��HdT�+1@|��~��"��c�}(�S5�����ڷ��>�n�\�7�� �HI�G��{���ú�SJ�'u���gJ�.а�����VZs�Ke�)�/�S�x�_�s�ׯ�~��c�pcL�ٺ�\�:���!��%�ʋQ�@ޯ(+�����V�<�����V���f#����귡Ǹ�l�nlX�l��lᴗ�Ƿ��BB�����{"X_��X�T/'����Q��DW) �O@��H�4�^�0`�h 
�^Gou�P�6�߾�@�9f�[ў��(Híp�&���xt2�b�>Nrņ�`�������m�k+"`h:�g��{����)^��w���w:
^B��?�0�M��K��0M���r����z#�)���ڢ
�z����c7@*a(�� ��K�A!Jȴ��x�W��w��M�}�ABѻKP�C�r�������*�{���5Ӂ�J������ی���"V��;?6^^.�$��;vgz��X�/I ƣ� ����Ԑ�f��q7|�|jRy.P��}[�{/r���(�p�];�ܓ6$�	q"gK3,<T�0����7�;0m�u��_�
�ȇ/",����N�l0�0:k����;q\Ee;��1cotɩ�L'���[��.I�8o��j�݀���#��� �h��i��@-���y�>K�}g�D}��Yʟ>\LZ��"��/�;T��ϊ.ERC��&r�M�-Z����O\���uAc�c��:�U�fNО �jɔ�W�P�~7��������++� {��gS�ѥ��s'S�hX7q�s�ѷc6D߲��(�뭇��A�Q`*�Ok^����.�����!O��2b����<�)��U��X��#����|��|��e�@k�C���ڏW�C��X�/���ΎM����`f'BB{{�Gg��]at��qk�.؉}��~pX��q�s��B�] M&��Zo��;B�[0�Z�\;�nDo�#���E4��T�Z!� zS5� (W����ݽ1�{s�
p������_���yQ���;�1Ҫ�fqM��3|��+y��c�fs������NMc&;On��_	B>��sc7�T�VJ/�5����zD��f[yw/I�����9dd}S]/1^�t��8������g��6?�1���8�b�?�2�Fp�l�V�$*JI?��SW>�@ݶ1^��~O���q~c�Px ��ʲR&HT�GN����vbS�8~�^��qBH�qr3Il�B(��"���޲��u�w#���mO�E�P��� �å)P ����׃�?VgR/�j����d��`�/����Fr.cC�3�d�V��~��}���/�8��=P��g�qQ��k`f���<�Fw�1@.������m���  �<��'y;#��k��.�L�����U̵�UضC�t�v�_/�j�XTG+�c���^4���ͮ8-��o�� ��ST�y7(i��̇r!�R ;A@�E$���w��W[)��^����9�f��Þc�,,~�߬G)�>h�yO����A���-+��D	ģC9�l�9��!���/�V�I�vq⦩��$ߥ_�ŕ�fT�-�R֔iJJ���M-lP�@�AF�M/IU�[/����ҡ����M4x�\U�x:_�&c��6�+	���VX-��<�厅A�����ֳm|&L}4h���0����ȿ�7@����.�~�0z��ɸ�-��}�#��S�k!D���U�A�G�^��$D{_���W���<Xm�=d_����YsYQHdx����v�&�<���1mX3�=r�'ԍ�������@��@�=,O�����`��l��&[��7��\�����+�����M��X��k������W#���ND�{��O��P����7&DO���p9�������M�"���$Cy�o�m�Rubw*�f����O�Rn����z�nY�-���&w9�A�3�r��_�<�gf��Ty�"�=n!�N�Q=��d�:2�����5[��9I���Z�&����h� į6�s�M�:`!v��� ��{Yr|v�#'�pq}�E
7��3�z��tE���^x	�L2�~�,���k��Z3Q�(�����->�,[�0���,��Ib�׭jq��yvb�,��
�rkX�r�x#���z���e�jKɉ��l>)Qd$��~�]�rp�	dd}�s4d#�Oe��`)A�@'��t��B%K��d��������,N���e����%��ϴ�O3(�~��Bm��ײ[������ʏ���5Y�x�J��=�9<��sk�h�9�)Sx5�7{�C�9�]�ő 'NS��O.�g�/Ц~F��i�2��%���Upv^C� ;���a�k�
��6C[����}���od^|=��m)_-G�[���ԍ��Y��� �7~Y�vNտ�mՀ��X���cW����
�L���Y����FR1���b��b�q+C�?k>�$q�������4��si�E'��g�t�q�:*��8/��vYEMU_ki]a19��6�JW�b0:���b��w�S����;�!٪�9�ا�$C��Y��1P��L
�� �fd�VI��7^!�t`pc���!�jf*������WjOS�7��|7���ķu��2�� }����qMg% 9���4BZ�
������+~SD������k51D�4��W���&Uo�Z�K�;U��4�^_�C��=%I�]���9��5�OO �N�X�A����y�y�[�=�B��E�'�|5���J����O�u
uN��l]\��Y�p�܆�~)�W���C����;g�?�d����Ӥ��o�1�����qۏM��ͣ!�mϵ?ݢ�c�e���յ
HT"��*�B���Q���FJ-�ӵ1�N��#��� fc�?�(�9��ΐ��2Z� �,αςxˍ���2̽E�|�0 ��D��`�1j�Z�y���Į���=O`�seU��ҫ�:`�O�^SZP� ��Ce~�W쵹��`���M�����M���\o	^�'u��#M��p��ó�%�?��W���3^�SL��~���Ϋza$�d��zv�ʪ�X��^g�*/��$� kv�#s��"{����Jѻ���I�Wº1�3�d����x�U�w��*.|��Bճ�����	��e�7"��G��q��wK��b^�y�g�1^9r3r�?����QϿ7���N���R��Ԕh(2w�\+�Μ�l>�OI��a�wY�?U�;�R4ZΝw����ү�;����^w~��j����ZS!5�;�k���Ǣ���&.�6�P6�+�
|���:ZY�w��&��zج����MT�mrn��Y����?7M����E�M�/��~K"~X��8�"mx������k*g��~�~+�����^*m�#��,�pc3x�抓?��\��(KC:2L�\�"ٗ�&	�x��_��'�5�͈�_�ըB�㊘l�W�wg�BܰI(����Z���t�;��I��~�W.�Jb r`���JQ��H��^#�����A�ǻ����%\�'ܾ�,��b�6U.��uD�ǝ�g,!�G:ӓ�/���.��se/11Zǃ�1Tw�F~uPy:��H��9�;m�{#�����w��cc���(�je9�����Ɋ(�~{bh��1�3,1�(�N��d�JV�#伎;��i��@�
��M��c�`9���8�ٌ�*�.m�}���I��*��P�~��q2gex����l���������C�\�!��x� Xp�� E�Sp����q�����Z9���&�hW�_7�.&.���`揁��&�/%,^|��"���Ûw8��!�Dԭ�Ж��Ϣ �f��:��w��/�Y�
0��>�%���@�F�W��|w0Sto��bd����U�Qb�������N���F{B�����4D�6�"�੶�ٓ�"�W�Z�m���b�޸�v挿��w�����E9@�n��9�͔�A[8
r��&��fdl��I�Z��Z�5�Z��jj��*{�ε��am�^��H<*�Ύ[-NT�F}]U#;���2� C����(�]�z�@�W�[��MPT$�9��1��
s��1�i����?���w�� �J^��Օ��9��۔�:����%�2���C��F�d~=����QF�FE'- ҉�2��&nw3(�����P,Ρ'��Z�v��%���/�F:!3�B���]^���l� -�002H)
�Fs�IՁ7�6���AA��ͥt�M&�z��g�L¶$�����σ��Y�m�I��%?�t�ߕ�זFG���'����Z1s�
Q׈s��Ÿz�n��+"�W�E*�uSN�1���S�>���X���gѬ2���_��=Y��τe"�W�����G�p�Y��]�����I)Nr�:S�(g'�7����I��v����)���y��E����nN�pZ��?�D)���kخ��p4:���TZ�'!�3)^s
���z�(��H�$;������4ڊ;mȁaͥDR3��a�\����yU�=4�	�_�;��I���EUb�����ԏ������#��p3�0ȹ��0��������O#-֠��`	V_Ԅ@Ehv =6�:�f��p�9W�ܑә���o�s���G"��ɨ[�_V�^�3���q�^ܜ���ZZ�RWzzB:o=���o��3��=��s�6r&[��	_J���vu%�_�!���x)3��,����Ah��J܊�L�)-��+�p���'�}i�:� ~��0Qd0u��<SK�_�Z��SA�[.������[�"y/K�����̷ii#�vӐ�e"V��U�!j�b�)���2]��~��=K�tE�����U_Nܗ����o ��_L"�jUkV�)����P�D1����=�_�	��$��Rm���<X[[���ʔ��9��'\�z���S����z|+CU�S�o~iS3��ia�O�p��V^��B��x]�(����)��ʏP���z�q��[���+�}D5#�v������Y�T;�K0��-'�2�l+��̻!P%)�oDP�{B��҂i���ɗ�"?Z*I����ň�u����E��:�-�@��C	�H�:�,���D�1��s%�y�l0�|��o��<�%����9w�y�B��I{z����J�o�[�<hg���"|Cq��Zr�f��~ZQ��� $�nĮ�� �m�������[$�MEQ�^��6?�}�o�I�aW�۰<T�`Q�ݭ����M�L��p�2����ͬ�	-ނ[7UQ�v�-��\nߔ;�5�W��a��`a�8�PL0���y���ֳb�5"3���(=崋uc��`qL�*�	Οͺl�p�Q�6*�́�lqq9)��JE�y���ZX�0
 =�xB�:$�ĝ�xyy8㰙/..�/&D��Ue��nS�{��O�Ue�/m
ѾW��ͳv0\�\d��?�4A&�^�k�9l���g��I�y�3φ�����CT,,,%�U�ԕ�n�>JV0�ݳ�n���e:�Eʽ�=���0X�_�f}��g�yߖ{9ݎ<v�]<�����Ł6�0ʌ��7v�W��Ύ
�㙆�+���F�@ddwǦ������tj����%�!ؗ����e�,�ɓ�W+�{��lx���ht/��J��~8�	�_�ۜ��60���{�2?n>q�7�w�wR>��D���?}�|D`�?o:�=����{A���9�t�յ�h����"�;9�%D4ז����Yu�?S|\2Y�Ũ]��y�ͻ�*1ۂ&)9������[��h��]��|9hf߱v�Mf�8�[����l�Լ2G��S�P���NEe�j���׀KVl�x�`i�#O�@ET�;-���L�f��֛2���3����l�B���v�m�_�	����y�'��o��}��P���&�Awy����qj~���M��������m�{�����׳G|{.|+Z��j�4��ןx��>\�Fx��A,:�#���>e��v"��n�FvW�ju)*��K��& ���`��S�k���zy���$Ņ��ԕ���ӱ��k��=!�h--~2x2�Z5'h����V�kgGO�|�M �t���X�d�,��Tu�����9+N�����c���,�����h��g�2�i�`	sc-�N}���\��=xk-bo��BY����*�M۵�j�uN �]y���o�В��L�����-�i�]U�/�`.�}K��gR�\�Yk���7_�����k�Zy2�X���04��.`o1��ϭ��.�.V�t㵌W�hQ���8\S,QA�*n�3�.�)���b�+`��Y`��A���~�ҫ�G���Q��ˋH�ڧ��Nf��\pw�v�őd]Մ&Z�Uqd�^'����t�^7��¼mg�q�������������ü�l���-<�F�/n��&�{�B�Ы����Ij[�����~F�7u�T���a�d��B����`N��4��6���'�oϴ>������A冐�~�<p���w �ͼ���,��zaŹ!#u� Pc��	:��n`�?�,��6]Q��F����^x�Z,׺Y�+�E��/��N+�;4��T��B�X�T �*���􌚨G��UDp�5f�7�|Q;s�<���a������W�$F�q��7�4�@7��" �h���*:�<wa�G���۶�k���=,؂Q�}�WL�hp������a0"���y�߭�r���7A���e:�5��$�~�����*��Z���=�K����(�g^����l����wD>�x�Y��l�6�k]��B�:��α��u�7�<�VF*63Mb���n��B�m�%i��f�BEz��	���� �ls>#X� �.q�Ր�)�ul�kʴH�s���Q�A�&H0��;���=:��m�pQ:�����^?t���޷�N<V�l^�k����EXٺ��;.�o��zYwƝ�0Ư���DK&
.{R�V0������b�ܳ�N�׻�{���b��v�G�Y�B7k����9���/���^�	��ԉ���os�����0����%��Q)�vF�/��wY�&��WlXu3�}8%a����ž,�?��uŹj�*�'lN�.�U�,zKֺ}y�ݵ�?��<(v[IjRc��a�+dY���	h]m f���m�g�^��?���-�Q�uL�yBb��޹���O/�����&#|�V��=�hb�ǡaK�g�ӎ�Cay�p�O��Mg�Zb2�n���}o��69h�����P�S�lFlk�򿾕�8ϯ�8�5W��d��-�<�U�����]t����"���yȨ�^�txx|�?�c��p���Fق���ך�Sކ`�E��:0O�����j<M�u%1)�"S_<P{7�O�\������q%�aI+��<A@�0q�ҧ��W��a1|}���C^z����uB9N2����Y�əq4Y�((�54�>�B��l��l�se8���L�x��+'RZ{�		�Fp-��|��/��?\*y|�A+̅��GQ{����"���'r{%�zX�6��#x�E�c��J.���@�[���
���}0��-7��T�Yj}-A�CNg�NX��샩�%U��X���ȣ���]�[;���x$/F�BP�?-��4������v�����5�y�C�nw�kg7�0� 8\%���	�+Q�W-B*������͙�a��G��ԛ��!���=_M�h|h���lĐ�=T��Z�ج~t��sJ��D.���S�_��:<��E��wO�����uU��0b/3���+�FN*��M@�_��|4��o�����l���2ȱ��\�}�kE��	Z_�k�{;��3ӿ2F���%���Q�C�n�/ևH�!�26�{������Sù�	a��j�w�T����Pi[q����45����i���Ј𝋑Y��2;v��moo/���s	ƖT�E*��r@\^�a��kF���b�K&������{	�o��}��ct��&�g�-��1=f����וUj����y��� ��u�	y�wp �(�/9�\R�������l��ԅ��X��B��k�Z'r�8��Ki)1��e�7��+���ѯ�>vh�����Ha��ϋ���$ߧ�ׁ�K�V���r��Uч���/(~ⴇw��Ŭ�����@0z������w��k_o;�&�<8�i�����?6H.�L�_���򪱴��e���M��?�Wr�S_f��� !K�	���㙁۲�,��,���ѢơL�'����e��Z��0��|�	�(���5�F����-��j
Paܵ����r�^�x��������=�U_�������y���M���ECx_��к�]鉼ԃD�e����o��W ���[�0��Z�I4X�b�WJ���t岱��}�%m5E	/�
��m,�� ��jֺM#tG��������&J�K����� �����ɵ!/uQU+�J�Û��l���S��O�<�I>Y�O��{�छ�<��O����=X�g�7;Sl$s��Zd)z� Ia��ݢ���=ڸreE�~x�Ǝ,��$Ҡ?R��q�}���1��=?�x��6,?
0#�h�lԸ��y��
��R=���8'i�Ǔ	�W�]��7Ҧ�Lr�t�\�|���;3.���1ki�E�F���-��O��J�*O)ahe�G�\-�,�6��51��S�Ŝ���f����9�b��D����ﲔ�~j�=���^��9i��f�~���}�a��K	`���	5!�����-�{��vU�R�*H��M#w��C�i��P�)i��ςDRqh��dm�R�7��'��rOk�����o��,��o�&���3���v�Z6�B"ǔ�F��I�/>S'�����n�a��Z�q�����|��x墅�ؙqx�叠�Rh*�NQm-&���eF���6��z0*�QO��;��[�f�����o�מ
zi|�|����1lƳ���|���[Oi<�4���v�GYd��'��'�:�xc�H���݅��*�^�iS���
��:�h���9$����wdN�Jg���Z�����Bx݃��Lm8�~c��v/<���X��O ��7nUī��\��$��*���ϲL�M���b+�Du������m6�Ҋ\v�^��s#��)�45&,��8�*T0���*N6Q�k�YM4����{T�����h
��\n��pJW=5���4��C����Q�����Pi��$Gǐ�n��nD:��F7��g|�����{;�9��9�:�h<��� ��z2ֽ�����������/��z4�� �&�۲�@�$���D���]4')�0����x�Ym7=�E�
p �.����/��^������8��WSߐQB�,ꛖF�D ������zM��b��/K���;>(W���N��-��������d>1s�R���lIŐ��.9�Zo�	)AHh���h��<�	�c4�TΤ�7�7z�����)>��z���[,�npN��O"�Q���T;l4�<�c���k|���|��Q�[)��QpDI��Gţ��%b�3�y��e@/��������;;g9:�k9�D5XƝ;D��@��5oi���
���^����:�6�r�QZ�܊����L��7 ���V�V�.�&]�{J�s�2$��ʊQ�n��8Q����ߗ��=���F���/%���Zjyw(h�p�PV� tƙ:�p-V��o�� �"t{�k՜��ly���T�n��y '�R���u��!�I��.��d@��hY;������ew��T��ڏ��
��Ga���������{4�I��׊Ȧ�}�(

hi�%�o��N�6q��ݻd��G����2��/�'�^K~�"E��LU�� _j|�X����$�<��K��߻S���6cUa;2�4�#��{~�$�Y�?B6��v�G˅���^h���!����7�&D���"�_qYK�}B�ҟ8Ű��I$Y�z3�W���~�1��4��	�$�M%���e>���8����{Kfw�LR��������ߝ_;��Sk�����'��ӳk'�1WlLQ��l��`"�O��m���RHY\Γ���ۼDZZ�9U�[�Tz��p:WO��ܸ]�<��7]N;?�����GA����x���(������H�y��Sx��nw�S�Ŏۈ�p!�C4I�(��q���Ɵ�	P��.� d�$1����B�����^j3�	��9K	Q��<�=:X��ځ����������.���֪]V�cum�ϋjG����Z-ٮ����Ӷ;�P�PiP�<S6"ȣ��(0J1Sˋ�=.Dpn�譡l�>ja���3��m2�dJnL�[h��G�yӯ0u����x�,H_�ҭ��;����x�);W^
�T:�H��~��%�~�U��.�h��Y���ɍ8�|���%_h�P0��a�Ƹ3��!�Ci��b��ۜ��.1��@�����4�]R*�o��$�H�T����p��*o�x�)��}`7�������㾵��6u����@���j\����d׏C��QZ�n�/VO�ev�t�h�b� �w�I�9����+����:�j�*�Ep@��4��N�	�7RL[�z��x���)��FQ�č�8�|�P��S,D��m��m���q��ɥ���䢞�X[���� @�mB:}��[���y���N.�/���P�����3���'v�qye�����щ%h��V00�Zu���g���_kC�̱���
��{ ��������n�����'��g]�M\[����O7J�CI�nF1;�rQ�U?��9�S�������4q�����^��B��dyy?S���G�t2�:(�	�+�[꘣�+7�FtfgHri��j��]m�[ I)��9>���aJ8�����B�b��@�
$�G*r��L�ˌJ��S����}?�0����sc퀧�ߣt� ["�L8Ե�`c� v�.�H��@6�5��m��v�}�����y&�8�d�}*S�=�7�1+7�2�p��?u�=��V������1����\���P7�RHvo�+I)��~%�|؅�M�%;M�Oqnɬ�}36g��׳�����a��+�ԫQal��a���$b �9ݻ���6�
�3bn��\��:�G}�m,�u��܏)L��bQph9����y��4�
����AR��yR�b�O�\���,���6�իv\�r�=�=y�/N��f$�z�]D۝U����D_�����sZ��E�M����0ϡFg�N�#�����ԏ�[��$��,���1���?*��U%��>���e2��7�����S>�6\n''|�c�l�A��z���w>�x�{6�s�dax#��V	� �����M?��FyQC*1 tb�Պl���h�<6Jz�im�񑟷y��%
��؍q��H֌�����Oٛ�vE)�6��"�\5 G����y�T�1�/9���J�2�!7�}���2��Ä&�qU�΀,��&IdT`�����Q9~�xXZ^'���ީJ��R�25MX,͎��1�:�c��~%�995��°���Li.�F���{���Tp|ݪXc�7�,8b�b�Ѕ�UȤ.�s5�!b0S�� Y�w�<2af���)�HPET9sP�5�7m~(o6�K�@�m�#Bû|*�RIQt�<)�|�Q�:P[�A�3C0�&~й��?�>��͵����U�%��w�f�i����-Q���<�=Be�{�_����:Z�m�*N�{F�����V�&*�/{Ѯp��)��M������ٺ~-g�����[�V�ǿ�� ��ڟ:��w���DU�ǻ�ǗY~b�.vr� ��	915[P��Ɨ۽R�Ao�I_�-�t�sQ��O�*o��������D��16ܶovVôԤ��Qy�%bN�8���y!غ[���ѽ��I�+���.9�_������qE�rA����?3�j<~�3DAe^zڳ��-|�W@�(YR��xu$Ő�"���.�z��[0!/t#lc_��F6
�2���r�~}��t��P_�ZB�r���s>��j?��c��WtD�
 �G��Y��peN��ii)�PA ��&�[�p���T�M�
�Q��^s��}`��H%�d���f|��F�:�ܩO�T�e��ٶm�N�h�.�F���v<��ll�V�k'ӭhDf�Z1P�aZtX�	���ǝX�'Ϣ�KQ�f����0Ƨ�ُX��ߩ��}�w���ƺ��!:�t	"��2�Zw�G�=~X�ܜ��j-��{wQ��Ȇ�"��תj�ܞ��|cm�9�Zz4���!��i����[AIH�Ц&2� dD�n�U�_̪�Irg&�3�H�Q�)f�=��?�L�̟��6��
���ȤDϞ �����8����Pp�N��T�椧w��d,�;B[g�s��#�5���V^�� �K]G����r������#�o�Qj�.y3�N���w�鐹z��S�� aV�R�_���b>�eG��������Ʀ�Zo��D���Z_�Hmb�k�39�[��Uv[�����

�K�&$��?ݭj�K��3z�����4sXUh��a�����-�k!J-��zQg��k1�p��`Y�ͰM|$at����XH� {g��%r�h{��FX�C����}����h�`�L���IJ���WJ�
M)��7s��̿[Z,���}�-1yg���S}��g�0 /�H�*�R�RȍH��'�ZU�9# ����X��'�b�ym�NA+�P�)���`��?�zh?���{��8�����Lwq��6�O��$n~X���|\[Ӕkn��=4�?$�\� 8iE�шY��ƄtcB��}6����%�����Xi�L�D�0�3�M�D/ϼ�F�-��f����b��.�7�\�

�N���3��&�D� �D����HBq�B/��S����3W�����+�s�}�]L����*B���Y�o���w���:E���Rk����l-B��O8H��H��Jpv�y=�&��S!��"*)��':��2����kW��	2p������c�[��m�yS��r��Iu�GO2�VC�h{K��Pip�p�t�J]ڱ����vr߼
�1{s�@�X�ԡ�����#��)�3d~s�B[9ݎb..�L&�<j�|؉0O�۫:#��Ol;Hx���(���j�_�ڪ�8��U�̃K:N����h�B�~uy0���w�nG��E�U���_����l'��(�X" �ұ ��k{�q���}�U�ᩛ��SSS��<����@i�:���μA��G��<E�ؘ/�sM"�����Tr-�i'L��?�'4��R�3�y�.���a�_y���6���&��JR�h��� gb�\����-:-���V��������r��eZ�#���0oT9��#�����ѵ[X �o�_|F9!a���|����<{��xĖ��䊹�����;@�@�LJ*��.�6Ń�)5b.o�-_�=���W�״�i�x:713e��Sѥ�X�5�s��1~�\R����5���n��E)4^o���;�c�:ZL.���r�ςikk�Ꭹ��i���V�c����trt�ˡ#����lua=�����%�"r�x��\Ѭ����u1����e-9��Cm��(侲e9�ޚ��O���4��<܎��@_�����k�#!;#ؘ�o%�^@�*��]&��KO<��8qi"'UY�zS>�d�u�la�_�����<8���׶v�x
	tM3�+(I�;sѶ�)Ô���P�@���{�]�(gYk����h�	dſ|�O�|g|I��s�����:06_'�_5Dqs�d<G������ʗtB��ۯ�Bt�̄s����.���,��͆'=$��Cj븗��b?�Ln�u�{�|�2��b�m���$���;85ϩ��'���PM��L5��I��?Ύv_K�w�m�]�7������#n}=e��p������6�"�F\���B#�"C���^��!K�SK��Pf�"�%7A��Mt��
�n���1���ƶv�=!Ƹ
��c7�W�X�yq.��M����Ìٯ}��3����i���Ѣ�z�XBؽ��|�?�������lA)��(I����vS(H�e�J�rL�y}>q7�VJ�-��1^�
G�-���V:,����
�iqs���|ԑ5��da9g)_��.#b{��4=��������{�	��6�ȅ�����D���(�3�"������223&�4�@HS�2�����Bv�M]Cչ	��Djs2�Z�s�]�Q9�j�9vFT	�<X�Ŷ�����0���c,S�A��T���72U�Oa^p'Ml:��������*�����Dp��pI�"i6�)e���@��˯���&��8�p4�^]5���xo�F���tp���\?|r���D���V�s}K����z�GP����~Ҝ�(��=��5���Z����<��/��g ���I6��h�s���כ�6ܲ�o�ݯ����qT>���C+�u%Y9���)�Q˛��=5u���E"���[P�_҄;52��F��>�:��!c <��*����hLK�>QE������;��y��W+~�
��O.<c�ݏ�wj�n-��{(����^ݷf��'c�ZBQ�T@���r{%m撥�MՓ��ذ�ھ�#��y.j�C��5�vA�b$���m~$�4K�T�>X@U��N��d��w�}n)��{��/�>���.��*%/$7y�)�{֛��#�D�r|�K���I����5݋�9�.qp� �է@�KzO�>-I�ܠ&�H����S�y�ܰ��!"@7_/�MMO���oPe-�]!0mZ��ir�6"3��X4�#/�AU�v��l�&PF�=}�9�=b��~�ϙ���LM.��ۣG��##�5�Տ�,T�� rh�)X���p�����5s���\�÷F�
;:���Q��2ܬ�열��~,� �v:g����\�>�ᠷ:��V/�O�p��"�yil�X�Y��Di�~�\�j6���&�R�Oyi������m!v�]�*;���0�Kq� P���[n��EV�Sc��b�ge��V�`1�r�	љ^V$K���#��f?�7`p�cI}��[:S(�%���1G!�D��%����j�����綧��Oq�H���1��m��~����Rh��d���p�{��Q�7��7��n�c�o�wdJ��Rmh�w3^�:�:���jF����)����P޶-7��P٣0��#踀���z�$���P��-f����\O�G0�#��JYA����]h���f�S7�Hi|���Y�>\�p�-N�����b�ddأ�d����2�A��:��/��vM^	>�Rj�b��Ge�e��u;m_���;�`�*�@�[<��3%�]Y)4N.����uz�#����ww=�XRKl~��6�q};��k���.��y�[���ΑG�=�7z}�=	�E��;w�CXd�r ]$����W�T���E˺3��}}�Ȇ$��n��Zͫ5Z����t��,�=#��sMaX�>drZ��~E��jp*j��
�Зu~6h�߷�[;�%&!y���QB�-�ɫ'8P����M�ҝe&U��MR[:���
�b�5����*QbO.`I~{�t�bY:�na�ǘ{�]}���J�U{��M�- 1R2����G��_�jA?���X��U��t`Wbh�v�S@��҃է�����nՒ'oH���nv�}w� &���g'r`��x��z�eN��}~�^�\?<Oq� �#���bgM�AAv��6s���I���]�'x�������R��!�(�W�*�"]�	S��8�~K�%��5y�GAMT��s�(f���͎�ܦ):���9�{���~�׮���[�G0s��G[%G[%�����់l��,�iYqW�+�p�#�g�1%��y�`�P$P�d�s�ģ�Wn��4-$��^�	4bE�>\b>�U��/�Mhhg[A:�o��0���hWz[�����*��9w�]���]������VÆ�Rj;Se���(�Lz��?���҉d�/8��(�&�j`�~`΋+����rnG�u���}���~衃i�>`X`��m6<��;���N��h�MmZ~�����Υ�h()O�]y3�rVo�p�C�	b�>I�z.f@=���ԩ���t2ep�*̐7ò�K��h�R+�\��[�ݝ���%��b�Ä�y������=����~�ط�����.!�C|���r\�x���zp�72`6���/~I6rJ�������&�i}����)��:�C�Qs�W��[I+�7�`�_1��A�?رJrn��.�{Zr���<����Hc�D���׻7�cUĝ	ɳ��͍�*0����w�U����rm=o�8���?���~s��,����}�;�W�6�s-�'�.A��!l��m�s�y�ؗ�L�7�l�\I�ѝ,w�kF�`o��mh��Ѷ5,R�x�D�wi���m�Z�=b�#6�v��j ����{k���$e���k��kV������B��ŁNL<��+$���D����1qWK3�V�,�L8�߅(��m�(�/`�IZ�P�ƙ����̒��I����8��v}Ӂ-�*��
8�9�٪�{"����nU�w�2ЍC<4GD�(���J�i��j��<J��o��ٙ5�@��.c4�_���v,x�~�����ۙ��R�����鹺�	�����	�tAH�P<I�u c!Z���D"�LYQhH����I��@+RZ2V��z���J�����蝚�ob�-w�T��8O�y���|��=a���͹��?��d?� �М�<({��F�_`��u���#��(�V��g-%�z������j�y�-�;
2Z�p�M������a^Ͼ���T:�3�����r;_���':�U��"iW�+N�ΉA��lƚƨ	�z� @M��Q����81h���_�ܣ
��y�Ϋ��1�`�>�� %q�Ƙ�����p���d�a˭�K��Ki�7ۣ�&=�5�jƒ�d	��wzS�����	�?Yv����z�E�f���0G�[x�H3���}���q�+��Zq�	U�*C���f<�{S�3�au�&�l&�⇒`/'�@�:���q�A���|�K	�H�D=4J���^PT�Y`��D�O���{}���of�Aj��*ڇb�ڹ<��������Gҝ��U�:��@�>������FLە���V�d����8��GKf6�5���<F5� eBN��;{rW s���4x&~/F�)b*N|���M���p� ?g�o�F���糮�J1ny��ȕ
�K�h4J��n}Hm��:��2���S^ac�!�{q�B��#��,;so�'Q� ���5B����`��/���������6��|#���2�՜
�;o
���|�[��xF���К��A:?�EI�������)�q��ũ���$W�~Ŭ���̐R.�$�:~�p~�\שa-N�[�7���;
�U���w�pU�O�7�H*`��9��Z�a#�v��D�6,u�v�i�f��y����y�[U�yUr����y�_��?�VɆ�Θw�]l4�0#�12|ii���k�l�p�!h�)a�m�^
tB#�Z搪�1��X'M���;ݘ���0����˞P�<X�Q;4G9������ N5�h̽�q�R�;Wr��~wT²����̅��q.�f5����b7��-O�)�x_�iMn�zA}��@�Hr����r�*c�3����f��sH��`�2(w��9�������;��ђa�f��u���F��<y��O�K���)�۴JW;�D�|}c.7�M�rn{�b8��,��x����;qI�?;U�&����l�H��MUu�<�E��Z�X�'<����	��I��Z�Y'�r��KmGA��f��8�|^�N��I�0a�Vޤ������u��3�7�P�'����yX}l?���g��[��X��}�t��b�����V�~"�P�AD�V�^N/�Y�(��;�ABۀ�'N�'*�oP�N:pT�W+	���sK�q*���D���Ò��1	��Z��@����ӡ4>ʔz��/
�^���k����|C��nM��8�7����N��?sZ�5����S77�:)#uw"�*�`wڼ�gb�tF}�b৤�Ů)W�Hf�f������.oy����sH�ٕ���*��DI�bRk�@(i\��^DZ�D#r���(_s�f�8Y�:WY�y���qi��A���/��'�6�s�QM!�3�A�vP�W}�AUN��MF���ت_�pQ%�+����|M��M�7��XVU��[)<"����BK�f�G���Ό�Y��w7��y=�5�=˨�p�P��P�|OuyЁ�m������-EW����&���z��9����9HpAV����a�aDޕG��:.s����TJ�ރ��c���Ԙ����� փG����h ���xKZ�.���s�qO�Ϲ�fN]7�#��R��@�J)�s�����:�qh
��:�������\��\�O5E��S2e9:cZ�������	U#h���3Q���T��A����A]�|������#��ű�bf�n������bI _��41���}V�� �_��>v}�K}�6��;kO8{|gDnp�q���Z!E\U͞3�uU��ϙh��)��@i��% A	q/���t��U]7"�#d.%�6Sn��VL1���0D9(m�$CR��s���?��l�u,N��m�=뺈�I���E����/���W�?��|$~�\f�k~va��Q��E
��(�JT����]�&�n�3�9��(#$1��
i�eH��Ǔ�n�v�9�5l���&W��|]0)���n�N>Zo���[lzZ%�./',>$�.F�׬������ߔ�&����s]��ư��tƀ\5�9�P�DK��i�V���R��\.筎M�kX�EV���&$��~3�B~,N�I�~©/�:c�1�6�h"�I�'vU����g��o����x@��tD�*�1I�a��w��R���UE�W*�I�X>Xn��M��PW�N�i�5�<BH�����ߋ�5�6�Ct�U�b'+	e=��d��eB5�,Ӭ�BڈUR��9�}gˇ��
^��`�d��l?��}�\�1�#���Al�q`�/�N�3���Ģ��6�8y@%�@����m#g��Cc��%�����˷������`Y/JI(�Q�f>6��	��͸Uc�\B�\�~p���|x�+���������D�S�(����k
�E�s~�������ZBCS9�@�K;�`���!�Q�_ID&���$n�4�
ۑ�`Ẃ׉��+6�d�͵%��7M���S���� o$?�EC�<�u���N�v�j<o
�V!�t��O�𑆰���Q�>�y.&71)Ϥ�BU!���=.u-�D��Jo������]� ���ݫe�M�;YI����h�܀�>�lZ�;���X�6c̈���f����yxr��aD$P�z�ʊ��&n���� ��*��Kf������/kA��~��j\�D��^���{���ԌwX�I�\��rF ,�:|��!�1Rٙ����~��Ap���o#�tڲ������߰U?��'����Y^�qI�P���'�2�	`���Ғ>�J*�F��-9�2j�dU��f3=�@t֍9�Ŵ�<�y$�p��jӖ�ܵ\��^g3Y|7B���i_���xJ��h�6����^P���iw�1@�Zs�d���P�͹�G�w��{H�9ʶ����%�M1���_���?�*n�o|� ��,/v�˯��r��\�qU3i5+�5ńo�[*��V�����������-	��)N���#��Ž�n�D��.f��z�<������ϔdIm�a�܄޴O��쫤����o�4qG�Q�J�P&erV��	ei`�&z���M֟9��I��(���f��Hdu�}[�0ź���>4Z%z�l�$bg��gjs@��Y-��ר�g�B	�^o���7.pO�4����@!ta�3�MSj��1�5��j�]�V<2k��:Ǥ��j�?ЌݐK�d.#%���m̃L#:ڕ������[�Iob��{��uP"�[;:~ �%lR��mtq4v^qл�-.a�Tn���d�5e{u�6v��
���|�g�z���\�i����S������ʣ�p���vr�$+wzr��p������r��WM�Y��]~M�-!ǐl���%�?(n�}&#l&���`!D��$�W��S��L��ލ���z���#�,�
<�M{���1�*�p�׏��s���i2<�M�j.�Պ��d�.<����K�̉�nY�Y@�4�BrTת�j�y�1�`ǣ�>�s�D,ICȶ�ф�
���|؆��߈���=Oڏ�]��ZE�K��j%��(~UA:H?94��p��0�We�&�8^�q�֮��� �Q`���%�T�U�$��rt\� ��������ee��]�c��*?˷��*ꎪ�H|
5ܭ�� �oѧ�'u��-�[��N��?p��?6��/��o�~���oG
���6������>׿9�#Pߐ� �Z3��ꥮ-
�Yݟp�@��6��-�/���y���zˏB����%I¹S�Qk��9R1Pp�x('���d{p��N ���=|�[p��l)/ے��K�r�I�{�X�m�H��[��ɼ=�P�M�<�����h����4RQ�\����SE��-'����7�tl �:VCx���s�0�o4���~Q�+.�(�u�h���+��2/����eP�7zʤ���:�y�C�x�ɾ��al�[�^q$>�+�$��ƳԎb�}Wo��^�&�#,yL7�|Q��1��>'�R���&��/d-��e��ݞS���;��ށ��Լ?�K�^p��Up��ņ���AՉFآ�L��7ZU�,�������=WU�&p)ɜ�p�	�V���cH>P2m�>�^{�P��.�}�{%�M��{ji?������tUx�]� ���	��:7��!��jIT=��0,[}��>�W|:L����1�)�˽%� Jx('ח@GI½������Z$���͛ܜJ��<JY�Π/º����@��ӑ� %�����Q�G]a�B��R�C���&��"�咑F�����딮kT_���D(��=��H~FE��� �5�5�lt&K�M��j��]=��M4��$�N<v��^�)����LG4�	��]5K���m��d�~��:�;D���u�W�Qȍ� 1=��xL\'��e�j>F3��|�&�Ξ����xm���(����H�'����*��v[N�X,���7����C��T{������T2ސ���D_D�ꃁ܏��}?|�6�M±��~�X��i�Y]يԂ�=��FN�]���s��R��R}B3��^�'�eJ=��n�����2��_Q[���S8�֓�%_H�{M��o%�2tAa�F�^�rP6c��h��> ��������7f��p�-�Hxc|�/Sb̢f>�|r�����:���x�|!��cK�]R��d�_KD�)K��r���/P���zGߓs�؄��ȇ݊l� �҄���@�çU�V��&e~�*Nk�3��ӝl�(�O�A����~��7>���~k�_���&����	��GX��1��-��Ĩ��R�F���O�I7k���)�ږV)'�evt1�{zi�Q<�{!VX�P�ӥ�J��{������iF���O���!�+���V�6tRh���P�!}Jo�8pr)��=�R��Fה����F=���j��5B�t*��|k~�-��-�\=%I�T�"B��'�s��wG�C������۳�.M]�n"���W� �dC�ħ6��͇}��W��\���+�,�lH�����d�v���|"ؒ���Ʃ��n'��*!������Mc�Kzѩ�"eҜ	!Z�KT�{<R|wWf�J�����@��{P��ygCХ�R�>��#���}�lA��l���p"G�;|���W��Ŋ�Q�[W���v��)�ݯ�L)�5��v��gB��d��]y�t���P(4n�\o�8�I��W�|� �9�������p ثӕ�{(87������d�2���.+�0Kq�)�r�|\]r�M}␘vH��q�[��&�"晐�SFq�>�/U)��@W��f?�H�H����(^l���T.{�S+�8K`���b��pr^�dW�lQ;�::<U�?�^ihH�<�@���0�U���R^�bB��M��v�=*^���'���Y�7������� ӭ�6����'G������_$�s��*�v�vs#+�iHm�����a7�X+��2E��-�P�[�����g�����-��e� ����=K����:c�V��r�͔���i���"�A�,۞n�]�f��X����uhd�{�[�#k�2�zD|�4��_�h"��YD˯��9B9]�(�.r�J�{÷6Mg��+�:Yo���3=��z�N��$��2s�0B'O�9[��������%ȁ����*�覦T�̳�?9~�l&�C�0}%Y�C�_��e��<���qgn�δ�O�W�q[oV�$|�1܎��l�H�pa*1^�.}'�&f9�l�eM���
�R^4ԏ�U�.m�3��˫&a�?��Ix�*<��FX�����d�a�.Ȓ;�\�N*�+},0�JGC `{�u�2
gt�[��	��Z��+�T������[����&��@7A;���<P,P�3�ٞ��U=M2� ;V�B�	EK;���n�V��+�C�J;�Y�0� ���$w��"4��g���R����/-Mb�z*������/}Te|ޒr��pVw`"��H��@�%�Z�W����"�Zuז��aOY�:�9u�J��ih(b3��jo���E�ڽm�J
�o���e���b�d�'U�4t���:�U~D�I#�<��MjG��������A�~#-D:(�L�ԾW��ۿn�k�dy��X�j���;EQ�P��/��U�ē�6vŚ��a�^(����)�
�%��A�zm��q�)}�3bF<r��y�9*�����W�6�M��߆$.�*�k_"��"1�MeH8AcOy�BQ�FF�����|�3�bh?`�-[Ce��� ̎T؜˵��Vy��$X��;���3ᇗ�-6�Yw��2�ѓ*�����>�:��)�^	��bs��)4����<uOG8�������/���v�h2�M5��&��7�N��S)l��4�{m���ԣ���]觖3j�� ��s����/���@C�����2�(��n���BC�_[/�M����Z�J��in*% �+�'
��̪'��q{W��,�J~ji:_4zR۟�Jͽ�m�Z��X�QW��JҖ9��d/�u7��u���hj�P�D�l��Iv!$����T����E]̸��/�����2�#�^m2o�?U�q����Zn��=z.���*dODW���;hZ�&�S�H^8?ޔw�-z�$��I�._-/����	<[��'��<�c�e1 ���ͥ0+���<`��0ܖ�U9���б�Ƌ� ���CA�Ï~`��\�f��P �w�'1������ڙ'���w��|�۷���S�A�Φ��|U�e%a2]������hB�w����0����ҹ�^4�*=!��|v�8�k]V$��3��W�$��w9I�x��D�&L�Cl�T갯%e@R�+�����C���y�n�ԌO�h5�s�扶ӳB5�d%3$��8;��M��;�=�x\�+;QR���-�ܜ/˜_�a��\���d�b���%Yo��Qb�q7�Ia䨰Ƅ/N��t6*y���}%8��S�<M][[��&�<�/�Yr.���t4,��uS�>%d�~x����ji��@��������{���՛t�&�C�Ŝ#j��m��h����;�~����'�^\�ݲ&���o��-2C��2�I�Yg�hn����]D��@T�Mp1>��}��#��OĩW%���e*޹���]m�+���T&v@�^0/���]ﲬ��ut�[hN<H㇉��Сd�>�%�՛��i#�_<+ /����Y����B�n�[������}���sz=\�W:ϓy5�$�%��U8���%��Ť������U���k�(��j�ݿ��E���Z���HU�j`�����:|# =5.x��B��.��Sy����l�z��H`�#��b=��x��"DQ��#�Z��s���������8y���[<4>R>��VF0�<Q ws���M�ο��;��k�~���7M�7��T���kΫ���w<����:2�E䧼�h������p����Hź#9��`�vO��P��+�i����p?b��(�`�Em���n(Ky���\�u��ݬ����a� pD�	�՚��'���K��� �}%��r٩:s��e�9��*��9y٣C`<$����*)`n���6i��c��gc�:���_Ȏ��JP%6����[o̗��z����'Z�<(�P���Up��U-�h,�t2�[�~��!�7�Oq��M
���#�@��N�k@}��9�X���
���k�y8�AJ�ʙ՟��óю8���\�}���L]>a{l��^��n����d����Fz`/��ma9��4�?6��A�X�f�B�y�B)��WU,�E����P��6q��|�~_�f�����m�Z��A�Py$�����8˯,*}� :��Yk=J��ҍ��g�����56?׮+�P�����	�~�AȄ��@$]`	���P������-����{"��?�G�i�����Y��ʉ��>JxW[�c�#z�+R�]Ft��\�ͯj��|ZU+ːoO��'*b��}�3������5d�����+���^
�d6cTܪ�8ּ
(,`�		럯� F@Ԫ�,H��hmE���ߺ)#��a+�ǭ�\KZ急�l�����ߏ<��l�M��tՋv��ti�d�(J5��g����t��oy�2��[���^Nh�n��w�>��{�i��+�rDժj��q���j�7t��7�b��-�c�ڧ~
dWV[�_/���sa�����y�ގ� )Q{��*k��q�H�n]s��-R���-��D�x_4�����%��o�t�NS�������`o���;��U �>z,I�J*?�Y�G�W�i�zኺk����Xp�*_C�����b�����	���*��K7"7��f{F��^bI��UI� ��\��S�׍A!�ԉ�!� #GD`�5}�w�L׬ڣ�sy3��� =��o���a���,Io��[� �҉�_A�������T�#�'���z����Aav����SVlM�z��� ^yϿ5��D�V��D�I}?��K����oDu�=ءd����r$�\� 59�(߶T*J��fO��W.�
J��.t҅���У$�1��_����<n��~EC�4��FQ�W=�pzz��j̺>��nK�U!��%��Y�Ω��8�%���˚;l�\�T�>U��H
uÇ���#���É�^?~�y[Ki�WA��Pw�i����f�t C����lF�x�ߞ���h�O�՝���Uo��u�V(Rܡ���C���ŭXq�]�;w�����z��ߝ�g2������k��J�׈r�|{�"��쏞��o��/S�Ѿ�䛊��X���U����A�Po��Y���5H��2%V��3z�B$�l)�����I��;����k��j5�iS�Ǵ�.�ji�j9��▰W�o�:Yk�W:֥n�:X��H;�B�ۈEz���E��&�k5}ҕ"�H<#;��(a�����ޖ�&�D8�6G��9;|_�f�k�_��kS7@$�T k�Hv���t�`�8��w�]�:7쮁a�[����J����\m��r'O�w.�k�Ȩ�P�xՅ�ޫ�����Cwl�~�� m$x�����BHf�e�����:րi��qO����Oz����њq喾�=}���R���5r��#�8�^��e֪��S�Y`�1=��	yeeZZ�9ƹqM�4u��[0�K|�����(��[�<]�(���I�M�G���ѿS�����^�【�g����Ɗ3�Q���]��ߦ7�7��g��l�D-�-��1� t.Z',��2��Պf���/a��ǰ���N9�"4P-��3j�l�v��﷗�j�5�:дE@�Q�?4P_Rx<�>v�����BƸ��L�c�)=x4�$��H�[#����
�g�l���)� �/��{x�Ң;�-Io��q���ז{��v��f�g���1�[��	,�b�@�y����p�E�GR�uV��z|v�ldg�����w�6��P�u��Ϲ�����Zk����ǐ5i��q�=j�^/p��	i>_
���a'�ka��߮aM�?��>�+��d��R��`鮪��6g�;������Xp���|HCwU����c��Lq�ٯ�O�ܛ�6����Չ�T�Ld�YMn��Wޘ�q��r����_��%���<���"hwp��Q�(��BO�_̌}��makh���QTU�c��*T�<������&����LS�KmP<C���=..G���ݮI��L��acC��a�L��f�e�H��XoO[����Ewi����a��~�y �R^��.��b3^��u��@=���_��߆�@��3G�x�)C�d�;<�67�`�����ef[I��6_�X�8��?̖��/���v���.���i�FV�1�0���H�p#D���'xP$�e~s� Yش^���ϻ��_�:����]�1���D�+dx��]����rU3����A%}`��F�u�ju]2P�1�V�ߩX�4�@����������ҝtg�c�,+��N��A�JQ�Z�*�["���u���JUe�;�-#e��-����O����ڭ[H�I81 �,>}nEX#	D�����g��ae���o��Cr*�i�U�~`:���Ӑ1K��hRn�Ms���/�/v�8��,V_t۾"�f���Q�C5Eee�'K�q�h~��7aR�}[�E��#(SUA����5��;����I��UQ�qX1����y�I9�1����[���-~�{�!���7{G�`�1r�^��eD��Ɨf���e�}�J���ʍ�~ͬ�Y�G�o�:-���Ս��6u�lB����3��\1�*sЕ[�-*�����[����_w9��q�{V��^]�xrgC���?p/I�4�Y�����'�,Ci\S�>�%�~���+8q���F���#��#}��so��NH��9O[pD�ƭb㔛��El�(Q�ߜ��f_�)ů-̃3�UȪ916�k�\w@55�/ŪX%�/�L�a�tU.gzx��R7�dɞ',xzl�m_�I��s;���b���U|�[d[�'�6������*8i�:��%�~?�)0l��c�Kog�E5�3i���":�ٴ�d�"�m�ڄ�<ԍc���I�ros��j(6��$���z�����1wl�~��a�j��%l� j�y�m>؏�*2�'�[��~&i��h��y�@��Sӝ~�h���>�W�<�����M[(0�g5�=���6���BX��(ٷ���	�^�o�����I��6I��B϶���T�������vg���,+�,f�����U��y�`Iu��5���c	9�	�nݴ���(��q��M���x�ϙ�u����>`B� ����mUa���_-_xr&��)��eD�S��[&>
����|[��^0Ll�Kh��u�!��k���f玜���(3�q'o!F��Ʒ�'�c��_�t�UK)̙����C����|�»W(�B��u3��V >�	�8d�{	.�U�,Tj���y~��g4�~DJ��'�aȵd�E�N`*v]&ᔙ9�,��U͔g���2'��8�|C�gR׶������ LY2��v��X�N@@Pm9G�y9D�nL�+	S+�T{0.�E�~ ����2ôy=����D^'V`����.C)р���Yy�ƴ��H�T�H��-:=�nɌ�n]a/�X$B'~K��d��@N�cϪP�_���z����#�߁C,�XϷ����zneIFb�1����7�����}#��I ��i�'�*��U��!a���u��f������ij��mhZ���7��yI��dx�&."t$�H�H�� Բ�9�m�7�,�k�TL
]!��)�F:R
Y�2�9�B�/�����+�u���Aqyy_$�:t�#��_�+���ő��r�LUm������L�	��p����Svpȟ=�SH!b�GD*�[�|#���ض/����\Xx淳Cw�ϿYƃ��u߳�����W\tp�))�5�>���;m�-�W��6�zC���y�_����0����N�Vs�>c����AFH�!��9��Cy�x�������ۢ�WT׋��@�Z���h�vaF�W�?Zo�ݮ~�Yj��.��8���"7]c_�k��V�=!�>!�o@<j�9�آ�1F#���c�x�����8�f�8�ư7�GQ�G����� ��Tr��q����x/F�8t��Vy���*��k�;Nz����w�p��\bfcM�Sko�U��n�V7����J�jVv�pt�?�)ָD���n�\�o\/-���:+j�N-��J5��w)�:��L�W�-���I�,:��k�e�Qi��c�6�K`
�΅�b/g����UA���Qwy����C�d�^i��~-L�t�nX�H�T>��3~p�.�_b�mŸ@"d��п�Nwx$���5�����ǃQIP�������=�of{f���@a��RR���b��c#�\� � Qj�X�	Lt��o�LI��!�N�ZTy�]�s#�'zpQ��'����Ᏹ�[v������[�ܟ����?T��l5Z���'|��Ϯ��ȴGH<�߫W�E&&�L��ftv�i��*�F`:QC?�X��i�Iۯ���J� [jZ��y����VUw��� l�r���8�c��͆6�<�8"tы������̋�:���ҒB��쾔��1��쯟�|#~_�O�����8zGB��~u ���,��N�<oH��fk�|j�3��a{��ß|xu2�� �U��.���[�
���J�8�~�|�C?c����z],&:��_���?Egyi�շ�HS�c�QclW��y���4��Ђ�O�s�Ǐ�_�ҫ � ����`��	]�#�+�*�h��Oc�V-������ m1���5��ZӦ�<,��m`��r}t4�/<.�W��õBN���T��T�����d���:���F�蟧�'OHl1*QH����\h�Oa��U�����Bv&6���Q���q���(�2���@}���Ϩ��w�ͫ���x�끫��:��8Z��������Iw�/A鍺���,��X�L-�!J7A�t��p����1�1���E!ť��,�a�M����h�� aJcJB�Ll:u���5���Z���@̖�9�A�Z��Vq6>\�ff�v8St%]A��}X�k��78$�2�Q`*H� �n#&X�̹����O:��&���,��Qeyb(��ě��N�ھy'w��Fd�J�HOYy���_]���`O__�7�7���?�ؔcV��~'���6]$Wգ/+1#���Y���N�YII6�bΎT��������caa�����T�j�|VU���{��>��e��5�ڧ��}6�##uV 41{�0abW��������� �rE�()ޱ���1��{�����T�������v둈����@���rE�#�m��Λ�pm�qsjb�p����̡�`gb@P�DA� ���*k��E���vo�	=���Z_������"4m����Y�:&��i��|�m�%}�*�a�$�;��_1��ly����)���5Asȣ���臒�(	��e=��D��'@{@���N��m�A�O�]g2��[�T�m�`'�Ev^۶o�D�M��l<��Mf�ps+\��T�u��ؖ팊�rlD�^�;�"H�:�#ۈI�3F��)���rJ@�O+Z{D�������O;|��y������/zM(��֯�0��$(V�7}��h�ЫW̦���D���>���̪��Z7qW���H�Z�(ԁ�MN���㡡�X3K70�݇��������
�t͇���r-Dy�'FH�1��Șa;�[F
��ó�{5�xM/�"��:��a�tv��r�]�-
�#�q-#|��
��F�Β�\���*j7�=r�G�$!E��C�i��Lp�Ӡ�	h�[s�+ ���֢Lh�8Q��A���(G���Ä�G��R��,$;����3v|V{#_Y0�t;�-ꟃj�=��V������Տ�>��(��$1����!M��2r���i��MC>���\�Ș�<}R�-)�˶�P_�Z��	&�^,n���>��H7�I�p����:�j�Ս��������%�;�H
�̱GCJ�\M����1�����YQr!�߽MyY|�{��)�0���� ������C̱-'�JH��B�"׷e�v�FPL����(}�:%A�R"�_n���5T7���	�{�J�VH`��ǎ�`�.YNg�Hlo�j�)�b��5��w����@�w���S( ��kA�Ί�Ts����x��8�P��v찵l�� ����gO�I_ǈg�:(�Y �[���������`lO��<.3��76��9D�5���Y�����V=���_�|��n+v�.���Ș�~)U����g�5o�J}�"%ƻ�z%#��?Q�D�6���8 �U߇l���(��_H_�sW4��vfr �bE����2��Y�0:�=j|�R:�'sPs������nL����"�G6%�_U���@	!��3�M.-�;|?�����.�w+?I��N�*|�j:�q�0�2}W6�>�x��@vGvf~Rh��Q�����,1��`!b,[ws�R�W���w_vW4�r8��'���|��HUZ?�q��G8���������C|$"Bh�g�˓�Ƨ�eN_.�<�Ľ�%�#�t�^���]�c!fh�B��-d�~g�|�m�!� F����jϖ�"���~���Q
��[F��l��}����;��ng�ʐ��x!�6��s��(���@@�{dz�F�D�Xp8�CU�F��kd4_����9����U�ݓ���U٬�>���ɏf���k��o���%`����/�!���G�b�p�m�+#���{����!�8I��-ɤ�=�&sL2$5&*;��2�rdf9@��s
��Lo"P~W�J99�Q%�x:�s�O^��_ڳ���9|9��D����_��<�6�9D�u}�����*��	��vMpH�ϵ��J�b��m���7H��9�
���|��;eF�.��=c-�z�=�~\��a�E=��5�6p�,�ujz��X9dEl@�	֪mE�bj(ƶn��d��T��Lw?���	�j��/�A��@�[s������8|��?�K=�0��!+P�c�#�?Q���7�}�G��e|&_�\.k�ި'�Q41�tnmi�%�X�׺ :>�~g:ml�/;C��mD1M�`��O7��l����
f�^(q�2�~=��8�-3�;��d}V\П����t��Y)~ƿ;�4��~Mm����d��Ζ ������($2�w��{s��XMt���\������$pV�d��?d��0�n�+��������h~��dw�L�\j���2��6k�����J^Ȣ�g���Am����9���ȁ0C ��5�AYmA��Ω��ʎ����6�\3�� ��b���%�.���\�mG�R��)ύ ����S���j��zY�����jY�:����Wh�K�j��H�fw�í�>�3��.�¢�ĩ ��lJ�F��P(�h�cP��`R���"��(Ivh]�N�vs�D�9�6�8׽�t��e��(1�M��
-`2��*�kNSh;���(�#E��nm��`1�p�ЏͫW(�`Hv�6��:? �HT[� ��e��b��)��i[���4q��-6B��)�˖�j�+PZ^�����2C�-���̘���=�>���Ft�����k�6�`d��sb׬�Aa/�Z�2�K����oKO�\�al��f���	���2�9�8�bЄ��v�1����I�� �W^ߥL2~Mۋ��}�GgI���bI♖��-3�n����n�gffd�[[r�gH-�>.o��uR㻙Xm̆n�籓+��V�:�I\��^�Իo-S����>I}�� �N�z�|����?�QZ���ME�]Z�o>�8�T�AF8R�d_ɜ]X����Ĕ�(~#B�P�5�l�`���\B$�sx��M@���_�ְ�w�S��Yg0U!����*������3���w8	��66�a�~�y�"AH���O�kPz��#u�a��3:{��/�=��}���hQ�u�P����yQ� O�;��p�n���n�L�'oi#{�o�ĭ��`�m'���MD�
纟P �{��MKӞA��6܌�0�_�d����4�~'E��j�����?��:�%C͊��ј�1��߶�*:���N��ɀ��nͣm뙨���9�I�	��8��$8��}^��u����@��,F���M��HĬ�`Ez�D�s���W|;E���+3(�bN@ �%N/tB��L�W֍��U��}����ַP�w��0��$�c�GW��n"(��AĬ��㸰>M:��Y"'��>���Fn�"��e��>�X�?�P̓�����J�V�����Y�\A�'�˝���N��/�1
:���\Є�~�����B��sZ퇿��<_�e�i	
�WT�{I�9�>��,�l��p��yB�>6����{)L��T��$�2��q�ֱ�;'�l�;��u3��e��5<�øl?�[_���
��v!�h��ѡ�^RU��a.fT�r��L��w>/�q`��DL8v�Kx��/
���� ��|����r�߄�)΢[��4p�ɥ�{|���%)��?j��~�]��K�^ƕP;�r�5t��3[WT� ���-���b���łd�ρV`k���K�L\ǿ9� Uk�Jɘ�"����w�_�r��Z���_��"���}�����A�w_@A�n�c/^5J��5��(�(����������Cu�w8"wx=�-��ۜ�ؑ��T;B��_8��a��&�Y؈�6c��UGM�/|��M�\��<��a"ɒ TcÝ݆As���l$��]_:���)�R.&$e7�V��O�-I#�������?�9OΫy��BV_g���$O;
�k��|Ujr�)"�OY����T� �3>�v_��Jky�^w�ܯ�d���t244|��Jv(7����X�/n��ao���%�
�/=�U`�&a� ��EN���Z3�L�����V�f�I�RM_�{����ĕ2��\�g{%In<K�[�T����u�w��ԍj�ܫ��f�k�b̯��s�'d�]ɔ~��zb����9� �JI!1�5{d�Ϋ;��L�Xq6779������g<e��8�8�-��|��UX��٬�i7��w��n��j�}|�~�\��MD�n����K2�>�2��^h�/��o���U���:�� �a���ѿM����	�-{���Q�;��Sm��	�,�2570��5�t4�Z����e�$��Y%��(~Ta�U��l�Y�t-�+$���&�8����:h!���^����R��^�֝��ļ����[2�[��z-x�ˎ���3����
��ZΌ.���I�lT(���?�-�a4{� "�_:�C�Hrn����:�����cƎLgv�~�21G��(�"�Mt�ԋ�TI�ʑkK������໎R)Pga�9�?K���n1��Qb�Q����p̯e/W�r�oq�Mrd0b�:P4�6�6Y�y;mdd��u����@�⋮;�M�׋���Y�EI ����wz�� ��̂��b��759���%���+�%0E���y+;�Lb�_�h�:�'n�YԐ3����8��l�ػ��i����,M�Y��ʼu	U�[����޴ �z��˱�qw �O��$˘%1��U�=Z���KyIs\���a�AT���q�K�U����O�����4E�@�GԆ�W7Y�Z�v�~�E��ь(�t ���\-v�h������?��oOX�� 2}d$+��	&^��S�
z���W%��TI6�ݹ�Ʈ��B��]4{��ۚ�������M_�u38��Q����^�X�NJ��_ĝǪrCm�����Xꠧ}'���
�����MnN����5�@�к�S.�1�`H��*B�����q�V��PR�p��NY�"Y�����%���p�"pG�ر�"����,o�$��|vz�?/��b�����S���-Be�4�}��C�l0�^\�O�˝�|(~:�<{�8�w��E�SQWJ��i��e����#�F����e�vg8S{H�L���垹�y�o[��גn���>X��_e�m�ǉ�E��+�e8�,�w�e���D����9�N�%���M�
�Xg��tG\&�����:���S���ZwJ��`V5������`���(O	|�SV>�n�Fuj����l�t+���gt���;#O���6���I)�Q��*=L��7Yt�L���������E���y%��?�;o�9!�N����ּMvL^�S����pӪ��7&XMD�G�0��#����7�J$����}5�^O+�V��R&�b���m,��\+�����(gV�<ɗ�q�O�h~[�?2���z�/t1�)��AeX�U=��q"7v�b�L��ܱk����}6ӷ�Ӧ�dP�s�C���J�%�xv�_��i_R��Պ�x� 4��������9O�rz�?YLa��F������힧[1=(wӇ̹�[��q�Xn�_���)���gq�E��,<�����zP[x�_���(~��#u�����K���?,��������o���鵓��rp;���di�6�uߖ�,��i��'z�_G!J�&Z�&� yO�c �-��C����O�����z���@�jd`0��f�'���&ЕK��L� �M!-�
Ǻ8x��б�lW�ۦ|���$}����`8>�Vv[/������o�a�)�j��ʐk�p��ݷ���UYYu٬�mi�s�!�i
I����NŒ3m�fn8����Lj�r���?�0��=�����0G�����v`&΅�.�~���g�"�n��M�`����WY�.\�I�ę�p�� e��v���վ�/iLQ_M����d�������b��%��U��oD���(�e�1�����oL���9��f�\�FV�`�pJa8�[�R��-��������!|"K]��*''��݈�R�a��STQiN|������p.���]q5�|�¶bv�Gn}�t��������z�f^����ǰ3�.K�H�g-���M
�'*e�*I�̃�����X����Ј*�(1�7~̲�*�0��;}H4fe�z��+۞`u�������z��2�d�b���}��b�;�Y�Ԑ��������vr6��%Ec�j�ülb�vGC����Ǫ�~G����ᇫ��m�i4�H�����&D�)w���e
�!"�H�Kϲ��%p�8��A��Wv�C	GC�w;�b��r'�h���h;�DزÎb)��Oϼ���:��K��<�������;m:�,A_�I�9���J"���}!�I�i��\c�a��G�eM`׹\��F�J<�4�c�O<����`B)g���.m�T)��� U��L����R(����a=���H��"��`�}`t�`a`�)<�F�}A��b��Q�dU�̳v�e��;urXڢ��9�ja�[���i냀�f�ՊLK �T�.EH��0�_��mg��M��Os����G`[�щ�%���@�A2�y�����M	zD�Ik?3$��vK�X�+ևx�J�o�,4�M�Al�y˙>�᧛M�t��T<E�C��tV�yl�gx�/4��(�� Dc�`"o������x�]�$n��Y�'\��ci�w).�,Q������m�4����H���UZ�1�gZS�'�L\�w��H:</���� �=�_h�R��ZJ�$���e�tM�y�b���{�"���k�M�@�_�t��,�S��oרC0��J;��H*��6���A�UW�<>��Xl��U��t�_ʐ������/�&��U��x4�Jo���L�OҀLl�E8u�	]y��v��"����O��Ih!h���R������!=ɫ���.T�����=K�
����E�!p�>��aY
��V͡����1�P����4?��� i�UB�lZ��8l<Y��Qt?!�^�<1���	}/b��r���M2�m*�k���F�X����-0j+d1"�ܴ���F"�k�;,�b��'�dZ��f�V��0T�Q�MD��JA#�#�&������m�wg�ղ7�8G�z������n��� &-Pd�^$+�c���q�W����1z���ҭ�Q/��.�?�`� B�G-��:���D7�*Y���1��RJ��V����ooS���?��$���o@�F���;����˽����������"�G6�w�p��Vվ�Z���HT��¯Y��iY0�%PBŁ��J��E�Fh�Y�T��D�����9��ߺ�n�z-�J��P��`�5��*I�i�<����A ���������eN=�%I��'��n�vi��Oլ�7�/M"l,��˶�5U��cʌi �ϗ�������K��ԇnQ�oB�LD�Cc(�%���i�'��L�A
���a=A�^A�z%W	�{\b����-��)�F��튫�y�y�ؤ�3�W
_�ϐ�˧e��3����K~}{�̗��F�6�Dr)z]�ێ���>�@`�V����I��E�
����[�/��Q��Nhq>s���c@L���[��e�WM��&�K5�,��5�8:f����L�Ze��D1H�Đ�VS��.oYh���m7a"츭;����-��2ޓ�Q ���hׯEgT�O4=�){C<���a	8/�$XTm������R��{��oU*=�w�~��-|��E�p/�1�%dE�~j�}�"X����@L���Z֒��$�)�����w�hT^��.a��:޾+�|3�\}E��J{zߕbnYe�����%����u�d�zY���n7>�a��M��u9،bs��������qe_�ؗ�6ܝ{�bc�X��y���,Q��5����~�*{j��+.�y:P�R�~�����4%�Xc*c���[�?�Fݛd��g�!]"���*
�y^�yDab��?&2ꆁ@ ~���6Y��%SŔ���Zj�j먗:��^k�LX���ΌFd&��(���"ȑ�&4�N�V//wn�X�6��"����p�2җ泽t2�F��D�-�N�R`y�h��C���&��B��J��\�p�a
Г�qJ']"�@Q?#Fܞ�y!ń9�#�ȣ�ܯr�g�`"���2b�6e�N�}eK��sU��*�HC�{\[`JN~�S�[����wR�2�e�I7�&���N�ֻr4�9�|~5��pꕼ���Ld��e����e=�X>ۤ�e�D�~�ڒש�3�>u�Y�iA�x���Ț��Pņ!�f������>��+�-�<-���~�C!�3ud�zLM-E�&��&m,a&�?~���ǭ2�K���sjx�P�Ƭ4�7l_�5#ܽ��}����`�xI@�7$1N=21w'���ik8�a?:��o��)t-s�M��D�F�x��Y�9U�ґ�c�G��*�]n���f����N=܀=�ݡׯut;B��*�:|4a�r�Jv���m�z��d���}M�)A|V��%�ޏ�.dD��(�$G{��C�0�����@c�ckfCm���j�,�q�ؕ��ODW������{�xyʱ��r�t�mVC�Y[[�>�["�����e�rDI�Lx>h�f)b$�
�䄸��P�P	H�Д춵-��JC�@���H��~C�Q�K�2��Y�N�� $�����t$NC�b��i������\����s���N����!4��\����]��K�b��C���;jK�9��e�0aYz٫�/b\
2�D����ܦ�V�	T5J{�d�����"�L{J� E��&�(��m
�I��H��ؑ��_K��5_,s7/���M�*i���-M��n��p�(�F��0f�sM��^���W`	���ܵ(��!f���\̜y}��Y���������.�M���H�y��Z��r���P�3^������×�c���|�U!$��DԄ�]C�����k�Q�T ![��܃H06����5m�v�?��?��4:��{ro''CĨ���_
� !�@�!h���D�*�b=��}���:���v�?��Aod����1�*���p�t�W��6��W�B}���]�Ug�#�@�X$�n{�B����'�����k��Q��L>hkJ��Ǜ]��eљ�.���?�ޗ�ds�:���,�V��|�cǻ@�0ٖjT��&�L��ɆQ5[������ F	8�:޲��~�"Ĳ�HEnFu7��%&�I� L�@�(M:��S����W#��A�h�W�b���M�$D��sM�["[i6f{�I�ZkLo���H}��`^�Ĳ<�#�M�h�b:Ҷ�WH+c湕@�L�Dn�K�m�٥�����|(����	=A�Ġؿ��_�k���DX��`�p��9��[S1�7�Ǳ�:֛�^�.�|Tu��센v	d���~��� �|�+�_|h0ڹM\t�!��Fex"����5HO�(�~;1`��M¢�A8��L\�y�����>)���yg�3Te�Cu���nЅ����ں{n���#�Թ��q��Î��h�=�>Ky�X&�h�W����cIb�ƻ�J� ��"���`8��m�(i.0A(�@j��������vͺ/�+8�0�$���a�M���3Qڪ��a��t�/1�i];W�iVy�jS�&����E1��*�NU�2����.�����|�E��,%$�6����X�^�G@L��sU����ep>�T��+ڊ��/�O����!f�J�Q�g��c�W�UVp��s�N�ׁ�|�(}��`q�����C,^�د�<ܫy��?�t}��7W㟲~^֢���{������>�8����DLR�*�ΟTs|���,{�w�Ͷ�TZ��]��@���q���F�!��h��^/��߽��k�c�$����[GfNS%��,��_���b�Zj�т�4�$�Q�����j��>��?��}͈�lDk��)����|~���0�uob:���.�������[���K��� l:���v=��mۃlN��2Z�k�>����d�v:��c��GU�t��j��]c��	�-7B�M7����?C���pl"�yK��QkM��jO�F�G� �'1b�=�I�8A(a	��O��to����yxZ��5n�o�h�����d��)P��+���|mu?<�Q]XJ��#��b��$�V!U%1k��	�ݻ��lL�`�3?�,ME=>>B����;�#��.����U?qG���c��/��������������Z.kr�*!��$WE�X�[��ۉ���qm�oa��n��[���']�I�AYϻTй��WR_�*	Whuw[�#`;�`:��Ѹ�'p��Lu�9����;&�
�x���F݈�����J����$9��]�$����Z�A^n�il�0~��0s�G5�i�ʻ�y�ϯw�k8�F &��[��n<��M9�s���cQ��(\��0-ڣ.o�9q��(7mh��,0,�!�KաM%�0�-���$���j�Xv�܋S֪��w�z]VQw�9�ʧ�U�p��O�U<]٘WR�w�4ef�'���4Zpo���J�?,c�]�gX��{��>��}#��T��7���
�LV B��%0V��?�j3!>�D���a�k_c�eHs?v�g�O�&��7�$z)�B;��T�������~����I��k��J�Iݎn ��xa���c`F������m+�A��|%\v�d��5F+R���w<���t�"���\�{>@]Җ�!p�\ť�
#oC@��f���3p��B��L�L��d��i'�l�J����ٝ�d�X��G��H��$PMr�69��,1`���Q  ��������oO��9�p��8z$�^l�:�}*K*��{�߷��?��6��ǿ2��:�~56�D�8t��[�N�b���a�2�9@��
��H�@4V�T���7����^�W$�̢t�&�����_�
1\���1��3�xt�Q?�D�W���r���p&(FO..&��9�z)�!>��0F�}uɺ?�?�o*E_�{���1;ܫq��cG,��,���R��`�XII9���a[���-泤eL�K$)$Yl�v�&�PR���*7G��W��F%`{��whr6T��q�0��T������e�+/�~M�D�Ғ�ko�eTb(�RM�ț䟿N��F�]2WK�d��]��3`l_{E�r	y�C�;L�p�����m��FT� -!�7�"�n�_��ַ�h�E^ΨX/|������2��������Q"豞��%:
�)��S�Q9����<�~�*Z���M�	6�=��_B�����͝�ۉ�4�/�Ҭ3WR������7�@��VE��?@��ܖKq��5Y�t�:�<	��h�F�0���&��?��XG���GT~��w���Y����w�?�~z��l�_M����ۏ{�O��^lbVBt_�;a����/�B]~�HG�>�	w7`"���ϭ:��[���j׭�+���׫���紋����3�4�������<���*�,`��_j�z�6m�u�,�q����
x���P�+m��r���<���*M`:���f��D���e!]/>h\���I��/vO��Y�������BvK)؎��Y�΂�C��M�]jgf^����W+:fM.Ic����p�a�_�[��8�}��  ��j#����7� I�[�*I����L"⣣#�#fU&��^dMB���L�*>�L��L��ZX)��N��|hjĎ����E�4?�C��.TO���ȘCm�-F�0Ϋ�)��]�C�6y<g>ĠPϷ�{l�MW��㠶2��w�$�Ƥ_�+�88��V4�V#Z�2��TʢT��U꒤6��a��7�8�� ���ˉ_5�$�!:=Zv�_w�T]KΉ���_	Ձ�hj�k	X��K.z�T<���;Ey��Ϭ�귍/o�ȡV��0���^���\V�f�krg�b��t���aR�����D��ڡf�.z����@���j*d�Y�h�@1QnBvs���HO�����s�+F~�Јj`����8�L?����@Щ +����#��+�dP�x���i��B[��IB��8�{���纞"�/G�ɵo��K>�1�i���P8�N����eͷ|�T���'�Ef�f�֎��|�7A ��7�����t�$���x�"U�:�#�������~��μ����&���}Q��g��;��*���$�VVP�aݝ��xz��<w>��ﶌ��Y���,����b�jCz���+���+B�q�tNU� ��z����]Ǧ�6��`F��d;��������xٗs���}�*i��W󥹸N���Fd2�f�D�F�B(��O{w/���{�!�vb��k �[�zW8�7��?b���u=,?�D=�8�V�K��l�K��}�] 9P�PIZ�8{h�y%F����^�UcZ��E�����瀚���i<�|܋3k�h��C͙>8Ѓ���PZh>�B:iu{�g�% ӈ�#�I�4�_}�����3���8��ҵ��ǫ(��E>a7Kd��N��i>��cX�r���}X�(Os�\��{���lH�zA�	;Z��L�šE_＝�Ma�;����n�ʦvx��o�űD�
w�i�Ǟ`ԁ�vw����}�JЁ�P�ջ�S�$����:��S��̪�����[ ����5���{qkq)�Pܡ�kJpww)Z�%-��ݝ�,����{�o�f�@&���=g�yvՇ��ً�ӡ�A>:.��\i-ч�������6�~�>�|#��B�u�{���e��u��~a[�������X�Kpmwi�P@�<�_=5]����T���%�Z%�h'a��+Sk{,�t�>��z21�q��5]D���B�/&v����g�D�|U7\R,�S������|���';��
�R"�{8 �z��4���z�~j��B�^�-ϊ�f����r�g+� :�NL鱸�G��h�q)ܳ���k,��m�C󂧺������mҏ�P�`Ņ�m @-�q�T;@k��P��B����u�O� ��/�#���%@ɻ:ߖ]+Y�b @��£�
Tc��Ƹ%́�q�r7�h?����e�:�dP�7ֵ�u���{��Ġ����:��OҤO�$}d���-GF��]�u���R@�W�����wZ��PB�3F�m�?$&��^�"=��* ��?��!�ġ� /�,T����:���&���:Ǜ���]� {Lç���@_�a���P[&�쨳IQ!iȸ��?=!��ݪ�eJ�n4����?J 'YY����_<Yxb�bvSu3��MW!�:�]�W��X�[VP�E=\��f\.(n�o�+iMdy��F����X(�a+ÑU_x˔oR�f2�EAj�%�<UH�Ǔ_!o��$;�����Zi~0����'� p��%0�X�'-2jo�_�&M~4�#ʢK�o���L҇#y׻�Kx1u-Ͻ��I��1�^n��mt���6�solQ^!���WS_+n$���T���|%6�)'�f�:b.!�q�2�ٰ/;>;��Z3S�~��3a���M�b�����xLV���#%���ZD\O6mmm�+;=�N͞�*�L�e��K�oc�a�Q&�]���n�����N�L#|����p��beh���)�7I봅��g�;^��QB�K�a=N��}�}c��n����!5[�>YMw$�@T)�~M��Ǔ��t{W%��&5<o\V�;?Op��˱lFC_^V����bk���)�o�Yi��������a�ҭ[���6�y]��VL@d~��4'�h��\���4 ˮ������f��k��*� (rI���ș�H[?4�%�k�.b�q��9@�,�$$Db�Ͷ����S���c���?���x�F�B�4hs��[��b��c��fA<lZe�]D�s� N%*����\��a���3��-2�O&x����F�bj��XbA�{�ի������G�c�}�O��(�J�F*��=�������^�q��毋����:j4�m�߼�/=����w�/1�w�
��7�J�`[��b�8݊���\v<pW1G�\�E��o�`�v�eA_����L[�h�8{�W�p��?�pt���d���@�3�'@a
�5���<��	1d6.F�&ԨMYt|��ס�5y��6��<�Kͣ������+mF��&$֖s�~�?Tl�u�͘ޅ�U��dj�ߨQ��v�T�{վ��;�`J[�;!3"nB@� ����E��f��U��G�AA!�j/�Ȍ�f�5-�g�n�"}Cң��7-�R�/?(��/UfgcUt��,V��}���?h��~y�����&�
�qC�2�4�9�~t&5.߹1�q�%ϨLY]�����$��p!�wc��Ǉ��+���U#pA���Ô{�2g�0(?U=����ވ��4x�[�t��<�s����v�,حLH�s<��vv���;�GM1�晭��	���#�0H_�Lj�ޖ}T��`S[�	�\���~�6���_8������R��	Q��f�Z��Q�/d��1����7�}�-�\/K���$
x�T�=���i��ϧ;�Y�y�e��򰆽f�W
M�q��;�_V?�'���q|S�F=9����X򾇺ެ�Pzi]����:)��~�_3�#�q�fX�5����� �U�k�����*�N͂�d�H�#����H���K��&�I�����+��W9N�W�
��ڻ$m��6
T�����t_�K�V;m˔��3OV�?�#�y��-	җ�c�-q>���8%[�5����հ5�񦕷���Ŧ�@���[�?0�呴T	���)�d[�E����NE��Yz9�_k(���m�^�*�@$�҃����s*K�ʁ��³M+K�Ll�R8�3�W�~��}�X�G��k|C��mAq��5���@)4�[L��U&�z��#F��aJ=ת�L��병O	:�[�8]�m��Ǹ��f;����ϪY�nN����ݵ������-)�H���������-;,2�\�w1�YJGG'7B�,g�[�_�{�D��YT�#���<飂��H�Wu�N������z�`kRO^(�`g�#��6� ��\o�]�ջ-
�k(Ǹ��=�-1H���\G~��*����+C�{�W3m
��#�\N��C��t�[�U�1<)$3�f����\��y%Ve�絫�N�H���OW�J�6��izf�x��V;o�/� ����|nl�7_+^׬��n����)�ՃW��8򥏂�ҍiE0��`#	�غ�^k��a7���	{��=n"�����nK/m0����k�^�!q��[7�)J�& /F����TF�ղ��p#n1_�Ga���h�2̃]�b�\)ac�m�Śh�Z����H�@���G�beת:��Շ�@U�)X�x�YUF*����Eh��B밶=���=�(�N�E�������L-!Td
c�5V͞Yg�3��@�|Ar����o�7����uy�����R(��^$1��K����~����˥�:R��EUv�ǉ!3Z�����9}��7�>�Z�FR��s��s�C)#���~�m闆{]Eq;�A1���z�;n�Q���b2���A�PV+���/�͏N.�Ə�o4�OJ0Q{�W�	��/6��]�5�C�t����,V�2�x88�1B��0}��Y���z���P;������Kp�w�D�_v0g<���})��Gv`�YvXT�HL����u�#��$'"؊K���C������=� s��?�;U��Vّ�|���m�����{y�~<�k�S��b�*��f��-`
Y!\�gq!������F���BTID��Q\3j�;���Ⲫ>���߆0�7X풞[=�7ܴ��!�zRsF����_өw�V|��Y����Zʂ��D��Vg�N�yHM�g�ʡ�#޺czԪ���*tg��'�_)�pQ\C=��K� ;�zъB��j`D��R�^D:E7r�R-q��K�}a��ՋA��q��vV`�<3��ǩ ۷��I��G�����b�����q�17�]��a�p���qlVW��/ED�x�ڴC�p�sn���2���`85��g�p�6ᴏ4; ��[��C.�w�v�
��Y�QtQD�T6���@�2��Cy�@�e��$JGn���)~�ἕ�=���p㸭�Iq����M1��E��CGۄ����M�g���蝡\ ��5"�}i<�R�9��[�nHĂH}���1���{���FiYe��a�M�Nf�CꎓC#&b��z�&ܡ��šZ�'|I��6����L\�Yd>L@|v���x+��xN��Ɩ��}�kOW�h��d�> �׿�ϸ<�4��8�=�'�n�|���	$`/��z*v��m���#��O.��a�E$$R�v(X�#i~tz��Z_�8pF�I�e��D�N�#G��{9�Nת�\s�&߄S�<��r�R�����}�`Z<�nò�2]���#��|>԰;Z�哮�T�R!~ʭ�'��x�Yԧ?2Ɋ��8^o`(�,hz����ƾ��w�NsF���,�7q៖cS�Y{���� :qoٟ�4<���8�D>Б�U�Q�����H��:g^R������"����)�3�r�wԙ�k�/��0�����0̮���g#팱�-�I�#�A��E-�C��xp�F|z�r�IBv�t� n'-���pc��&knYӊ-���)�4)�
7KM ��,nE�]�|���@(2�&��hH��p��x�O,��;�v3�}���|�e�G����Yr��?��n�}�br���C&b����\�����\H�	Uz���ӿa{5X�T�1�玮<��N!��\�ђ���P�;d`��G�J�Kj{�c6N=��C��`�,g�����B����[�B�f]�ն1�̑�z���˶&2��Q��!K�������⛿$�\�0������8��Ń����P{���I<��|R�"��R�� �^�>��
��qgnT��a������[Q���l>�6�� }��u{�.Ζ��m76����kvJ�;(�QWzg8� �""�F=���云���^ZQ~"K�/��	���d@���
�QGX_^e�`#1�BL5��_�ho��M��d6k�z�J�	&��N�o��eƭ���$���i�'�t캊,�D[�� �V�:*�T)J��%�uR����sP��j��-d\���t涞 �2;ӏ�������9�����u�Vv�^� ��}��R��Ŷ�����"�|��g�;V�9�ȧ?�+�N�r(agL�ǘ�A�+cO�\�R�h�����6Em�������c�K ��Γ�7�LKY(E��z�9�%�]~��G��j�w۫X���k嵺xc\\U���ى�����z��P�c��)b2�N�Z�zN�-u2��A�m�|���Mn�݈[��1����r� ������$���MFOꒄI���U��+NS�,0��N�ER�s<��4�5���G�)__�E�	C�>4(��e�!(�_�O�7�DG��$��>���|$4.�q�=�^�w�Wl��j�$���	�9�?xUk)�8�t���0Z��BwN����'�P�GOuc#vvۅB�M2���I���D�1����%qv�-$�&��ӝ�9�?�I�N{n�U��3T���ǈ?�&>^�d�En&�Ϗ�c�Fd	#k���덴Y�w.��A_m5C?�%@8U(ϐ�c%%:���ٰr<���9{�ЪSF���)6���<C�PΫ59�3��w�b�f",8�	�k�ǉ_�
#k�CaӤ�c�&�GP�{C%����������ڔ���쉚�ĦgR
�̽���h����P�7��a�,X��/f��'w(,�Q�_�
B�	����v���MY�j䘙�_�``��N$�Ig�2m�ǖ�@�B�)��|z%K}��70�?���H����9P^��zI��І#����{�#v���vE+���R�8z��sxff,\�dco��z9򧐷k7�&������Z�N�JWK���?�y����4���8�HC琚FԫD|3el����d`Ѫ��1���tw������R�����l��*�s��]L��� �'c�� ��y|M�%��B�Zߢ,w��%'�à\��߶%}�O*7H�J^_~� �@�x�^eɗB�	j ���A������{�{yn��L,N�X����F�{M�%$�k%\��kx��9��<[�>��5�8OW�,��k�cyܥ�տ�*i�����w�۷Ǟ���pO��G��DR6ז�~�����Jl����5t�"h�����=g�1�Ỳ��$�.�����WYMm��]�n{��_�ǅR��?��,Q_GbL��JO����]�+n���V]�L��r_����b�ŕ<f� ,!�dǏ<t'uV���ڡo1�ߕ8��ё���L����Żk'^�*����m�߾*D�c�3�
x1y8L�M��MH �E�=�l)Q�ż�Q��R�b�vL��(Y�d����7�T#֒:�h����9�8�[.*98ir,am
��4U)r�)1`�"HL�u���[k�K���%���w����o������Ff���,���ʻ��{�Pu*�d/��g_�n��@ه[�;��,�gC��K��"��Y�U�vu9F�ʵ�~t�4/��K�B!z�_i5/T�(�������U�G���(<[hÙ|�fw����Fh<ϿGv�]u�����Q3F���cЊ�������P~j4w�:�;`k1� �	��'�WY������(��C��n��f��t+�3����J�0��(,��C�rSe���s��.NV�/�/tU�>�P����禱�~ݱ�"�� Z��s�;�۰�f�|s�]����"�i=�J��5��@+�h���%�Z���ۦ:��}hPА��w��K%rj��,��2�(vjLzό�޶Z�lv_1�}�g���Yf����yߔ�6�Wt���!y��0*p�DV��w<��-�;�C�y��!�=;��4�䭞���&j�g�smޗ�r�zA���ףծ�BV��y��}�+r�l�9�ס����&2	2��*�;J7|ОJ�^�题�)�Ņ�����f�75�D�S��J��#��i\��8<o��0vO�b��D��a95d*Mj���Q8���/	ur2pm���o���;����bZq�K�Oʕ2�v
�;�}z��;y��@D#����z('����s�|��`��IR��z�k�m*��lTb����c^�?���K5�G����Q#��M���k�,�Ctt�0����K_�vTX��y-~�n uT��(Oȓ%Cn���{`�w�|HU�O�>�>�������l�uޑ���R�!ڤ�
�p[�*̋a�y��0���I**q	����ݪ�B��>]��J�Y&�\?̯��8x��ޫ���jH�Jcǳ���S��w���\t�%��Xv���	ؤ�Zk���h�� ��n��B�y-�l��G�R��fUH.�+���J:,�=�2A3��Q�y�Dag��;�a#	f��B�kn9�[L�fܝHڮ��6�Rn\����=����^]N��ON�z�	(���R�֚�x��>���m�� j��р�_:�����|ܹw�zTw��`d��٥�[�[�}p��bo�r�Ţ
A�� �_����+�{%��K�%I�>��z�'��>��H��L��vİ��O܀Y�]�� �]���d�~���A��uEԹI5�8o
ư�d3���@���X7̡F��!�s��3��#��[�h��p@����O$�"�zK�Y$�N&�A�%�[@�Pl*����1j�*V��ݿ�ݘ�b;�����;O�[�]�h�J�k������7�AT�:4b�uX%���<�,:�r����_���u��Ц.���+�ѳ��lq�T/��=����ߌ�꬚y�rȲ^�+�@�kUm;1;�?��4�
�G=�/Ub���i�I\�7��� �mx�
�O>Li}�A7Y�֕���V�z��x��.��$1i@J��#�S#�!�Ϳ�J�=����̹iJ҉e$�SI��_Bޒ����Wc�M��-Y�������?� [N�.Eu��B���}����3�[vl�7�ߞ���q��/��foVJ��q�|Up/�'�& ��nO�����{���2RF������\g���C�uB�����M�3���>3�|/��O�A˃��������B�>!������l��YA/f6�{�3t�k}P�}��x�n�G�/Șo�~�%�@���叇#lw����]��|�'�]�ln����p6�����a�3���,���8-�t������!�"���@TQ����Ԩ���uL���9R\D
�(i�ǣ�ܟj���Co�5ҁ��!,��l��������:���m�$�����v�r�,��������V+�hu����5�a�WY��&=ۖ!\����3��`�f�jX�Ϳ��9��w��H�T0�'9��*u�JX�z�^�����<��eХ�٫�مg�A���&x�4K�A�Ӽ�I��N%ۿ/��ĆS� �i��l�9=��
��gT\$��,m�G>����Li�Ù���՜hL�O���V�E~l�1�}�� _�i�B!�/��M�Ԇ'
�4�3�x]��C�evڲgdY8/MኞNu���f;7��d�k,%Ql��	����ӐA��ܲ�ё��4
����p:jQ���\=߼�c�8�q�Z\��	�;v�f��؀=W*ms�"�Z~�s�Uםro��*���1aeC���X�� ��E���&��sl�o|.�D�ʌi�5���v0�7�ϻ,�����.^�XyG�i�g?Ix�]�5��R�\<�:��ԃ��Z!�
\"|a�6TB��>�u..����|�,bS��A%�Zc>~`�.�j!�p0En��_�j�����,�:�w�w}�M�S}�D"�8�g2�	f��0Mz�T�s����b ��䫅��'f�?��
ِ�O�S3�Gm7��W��ߩ�� �G�O���dn�2�́ATF�W��ZחwH6y@���L�FUp�$�?K�~W6p ����P\SM����v�՜x[:��L-��8�2PW[���D˼(3���S�:� �3�R�y�l�9����1�����l����Jw}�ne�mS��	b��0Ŝ��܀D�.��T��w��c�,R#ng�VI37=��Dzi�gtʦ�`��$(���D���Q����A��68��i��-���9*ĵ_�ݩ�	~.�D���<`��A<�Z�[ً����S�{g�&~�c�Me��w��Fv>� a��7�4@lIi\\ ���X�SV��Ͷ�zN٣���,�̄6@��=e<ZVW�YF:%�AT��9�i�(�g�z$Fa�*M�qP{�\�@�$�j#��ô�oN>��IO��sk~,T샴?P���Z��k`<S��Yo�G����b�S�Yئ6MZ+�0=7���J�GYĹ���]g�y�
X��Vվ�]�4��j����m�t3����01(��|�~��d> ş�0�dp�;�OU��17�ă_��`���(��~���kμ��Ac)E�y�x�.}G?s�:-SEQ�`�_������Vө��Z���te������̝=�͋���8�����]����W�u{�ƻV����G����%f����2l��}�#ΣVbv9�󵈋;.�l9���E������%9NگC,:T���7�d^�w���k�*ͺ�#�5�����>�oLd��c4�'�՟J��D��|�$��4����̌V���+�F�B�4��q{�o���g���5悃ˋǩA�	�Dq���aF����b-c�b��/ʿ�p��g<J�\őe�9�C,���Kf#�������׎��d�h���E���suIh�X��|�pUlqqr�@�Y�A5��ʡ���T��I��{b��lC�S��m���g���.�c
�J�\�85�f�����q�h�iz
����]���L�W��/ҽ�ĘUsjN3�	 �E�j��v��ǲ�ҩ�-z����|�11n1�g?22���T�?j0�&!���L�fF
��8:���F$Y��������t�����੠���C�ړ1J�?���7=���Ό�L���9�$�"J�}ת��QD���ʻ8X��+���n�TW�r���0����:Cݺ�������P6F�hr�DU}Ԏ��b��k�Y�Z�*۟�r/A����}�	��[���c-���
7p �%+�aE:Ψi�_�s�I�r-��
h|�=�B�r,WƏ]d:5�8�����w׾�y����7r�����:�\�-�0�)��$��K����j�����<�)�t��<����<��y�M��Z� ���$���?I:bĚ~����^����.[��'�sq��=#�o�r�V|UV�ڤl-k���G�V�_�f�D�q���j�+W�蠮z��l=!&��L��@�?Q?��C�9K�����s��L����Y����<�Ǩ�wF���\y�f�(M媂՚K�B��3@�(=K�Ҝ���S��w�R"���uY���Aa��8�8�����*�a�d@+q����%lR>�	��������� l@���3!�B.�]6�Ԯ��eI3R�p���ޒޭ���  �9�x\N�H��x=�)�Hn��o����lc��u45C,���&��~��cqXw�z�zQ7h%�
��w�@C�Xo����7�~�C)y���Zq�]0�k�	l���������zN���Z�''��4r�$�\V�C�6���'����t��N'?���Y�+���C�ٌy'@�(�`�]����n�����$+T�`/PG���c��u9ca�^[CCc�0^�σ��韽X#�>c$c�Ȑ.�r�{u��c���b���|�ujTqMmMnELe:�@��p����i(Ԑ�9-�t��>YG�IJ*y�� ����K��"�6�(���!�IJn$�o����|�e��o]��ܟU>Hh����#�o9����g����un�vs�	i���C�i]���d��]�r�,v��~`f������u����G��|���
?'��k�=��������)�bHTI�. _OC�6E����Z뫵���4���}�,P=b�e�=:b��y* ��8�n�Щ3���s����x����yl��4������7_I 	[�2�����:mv����o|rm�����w�
�������Lv�c����	J�o��w.�)�w�=�5���Kk� )B�}�g������3Dw����
_��D5�q�)X q��H�َ؎z�2a�Ҍ����?�'��Scm��
�i��`�V)���}�lfOc�&$�5��a?e�h��!L+��MĿ7J���׻��ݐ�G�L=��2b��_���8��(9e ��b���f��ׂC[��0�r������v�M�X?�t2$_�y�"� You����s�\4��\���榿��8�fe���"�(�W��<=������ml�io�zI�9E4�"�|�	{��M��Az��1}�1��5��mơl�jv>�}�K��#�q�N���])�6�����D�� ?�����������=���EG����]�VX�p���*#ti�C����ON�N�}�٪���t�؜�`m���:٤���1�N�LT��a݇�e��s�IO�>���aQ��pC�-�w݌��-VS[����~+x[R� P���lix�&ix֦ř�B%5�l������e��cG~����z	����w�+���R�?� &��@s;X�w�1���c�
:7k��t/Me��Y����{�t�RQ���4np#6��ȳj��QU��xޢʆ�[�oa�qE{���_�M�O�P.�u3i����'���}b{G����b��n���Q|91�^W���I�I�����ާ}Dë8�'Q�J���Rd%!!�$�t���+"�ݎ�&��f#c������LV�*C��9�X�O�9���3�!�w����l7�bGW��:�R���y`�)����Q�]��$?���5>
r�����M��TN/8��+�����N��-���l��a��X1p�e�^G2E�5���t��ިT翇�-dh�v�K]���A���{�iǚћ��ޜ�0��c���ۭ���^�~��9���W&sC�ӎ�X��j pl�k��� 4��AO/�i�&�y&@S���	��� �	8be-��w�'Lԃ���M�~���H߲W4r�l̍������:����{ai,݋-�m{#-D��V	=�2	�Bv���M�_����M[	sCA�T�D��a>��A��}}�yI>����γ�%���S҂�i��	�z	�X���ςM)N���G��>�g�=ۜ���^E�h�oj.8����>�2˒������E>.P�|Ssh']�}����1�u"8r�����ʬ4M�4痃lam�tV�;�[�9���6橡����<�9�0��{�lfe��;����<ԥ\�&a�/����8��Ⱦqg�'\1Ps��`��)Fl�0-��&��;�$АE;B��΅$B�TY���#L�hiM1v,w�v][�{ ���6�Ö�B6����BV�PʅK�ۼ��W�sBH�'|ָQ�u]?��e���P��o���MZM�c�Ӥ��W;��E�xg�WI����r������Ɋ��Q�Y���))N��M���	"YB4�hi=a���JJ����O*��~���t����z�)d;��X�s ap_�U�UwG9+8����2߰c4�opru��D5���E���"���	`��ky�"��<ݴ�&����+:����\��ؐ��g��)�X949�����ڼ�IF�mWw
����N?�4�M��v�b���t�N����_��֭��W(4�z-#@����}���Q�Pt[�%��zڃ�8%ϵ^f�h����&��|:	[v�G�F�}���XG&.lI�0�R\G�f�{�}2�_�߾}�Y�3b<$A�2�p��H8wXi�˄d�9���N�K�~,ϻ$�mw�Q���~h�ӣ���-���N
tƴ�_^��������?���^���U�y�r{2���=�a���r��qO8�|����� ���a����o�!����7�J���{ay�T���Š�||W����F����4r�2�)�{־����"姯��:+���!���~ E��-�-�7Yr�ʧ���F����%9�ϵ��Ɏl%�B�ٷVu�ƽ1]��T�$R�Ĉ��m;|�/o��>�4���T�	z�|��RXX(�#�i�ьF��t���B���"�k���`��۱��u!ҕƳ����FP,��?���ܫu���.���|��+eJӈ��&�A���v���,i>=�e������O���i�Em*�^�hMV!�%�4g>;�!�x�*s$�Fȓ��[ʁ�bq�K�������� �UQ~�a��\L�$����~лSM��)g�R�����y�H�BX
��3|%�!���x\P����(Y*Wr���#8�xУ�#GKvc,KvRH=�J����(���J7
/���v�'����M�p���Dyp�sI����V�gQT��H�¨���ԣ��y�[�/:�h����	o7ܾS
S׋��b-�t{fQJ�"��W]&%v=a�U�2�ý�e�,3)�C�i��A��]�0^6�M���*�]�E��������;ڽ6���]���r6v��{9���Xh@�>�5���Jb̕7 a���J?ͮ,�%ē{���Q%�x�!�x��?G��*����{�Y�^�ՖJ�XpBg��f���pa@�D��9��RB�KE�V/��D�!(tJ��nQ;��
s1 ����-�B��+��#�8�p��6�"F������aQ��7�#{i�R�G<�ixa��{T$Β��J��"��0쳔H���y�y-��E���!	f�?�9ԓ9�����3}���󯔍�G��P(����q,}�p�
I���9�n#�N�]TdO��_�z�v->z+�k̔�ofTl�da(�UƉ���Hwc6$T��g�R���t����T�����ow����ߦ�*,���\����{��!��r��p�^�,.
����R�bk��� @�WL���:��Ǹz�鐷�Q�:�����7&91~9l��v���Umm���M�~(�� I�V�-�#V��B��䥖<�'n� ����NA����m~�J�0B���p���`}zRUmq�M�s2~a��8rUT�r�/�c�T"���k�<�l�R�]���y=��23k�aYGo:ƾ�TT�s��Ė�Q�/H����iV3U�ᘘ�f���1nbbAo�A�� Gz������W[������#1�V�� �gٔu�e����I=����2fm��8
a5�4d�����6 mR)��_[�:4��<�qI:�o���Jlb��uk�k[��0�J��4%�����?@nM;u��x�%砩�M�p�.bu�q-GS�r��������D�g��i���f��^z5������3��O��\��yb���w_�;�Aٷ���ӓи��`T��A��}���G�$�&���u;ݿ:1Z��2�`�?$+��C�f�_�H��4�'�)��"2�b� 3��`:y��R���;p�Se��q~L��%qۆ���w�&L5�1'J��n�u?z��]RTV���7K��]z�Fg�IoyQM��'*���?����Rȏs��n��U:�>�x���*Y��ъr.��2��g/�Ύ"�Hl��e�Zp{��@!_��sP['kI���q"~�c�꽥;fLV���4Q	�S�.E�wq_՗��߀�R��qY���8z{p����kc�#��ԋ8�lF�d��Ǫ}�FW7�O��m����-$����7��U���I9(@=K�����܀�&�0n�����s��t޹'J�A`U���l$[��<^:��)2Ǐ���~�A,A遁��I��p⩈"��4[��F���g3M]>���H����sf��6.�%z0�`���y�'��"E�B|��� �����@���{�/�@59!u��_��)�C�y.y���zY�xO|e�����P��+��	E������Q��C���%ũGtU, 0w[^^^dd�?��Ӷ/�)�l/#L�".)iF��@�vۗ}Ƈ-M"U��p6��x�g�;���̻ھW���o�^�� ���e�T�8V���I<����vjy��,��~�e��ߤ�	��a	��6c�u~r�v��>��j���$Sm[��D�<�h:�hnwf�l����+u���k3q����a۝�r�E�8�� " ���+z#��y��}t��drP`���^ ��|���p�ij���a(����~
�s�f]$Zf»��R�a?Gbe�m������d9�mb�7:�`	1{�
���ge?�q��T�en�;6"����H��A�ڹ�E�a��O��6�6%-�Z�q���m�ʼ�����5h�8
�C!���6}�~~/�_�=^	�πږGo���cWBs��g�}x㚥bGw�p�{�kG�ϰ{����#%��&xiCG�QZR�o<�4p�z�߷�fPDs4}����\��p�}V���!�2��q&!������c�51a�{�^<��\P~)�;Z�\��T�;�7"��J$�����A'�uԚ���w��+������ ��T���Z�o��6k���V�m��a�.���Oe��*Gv(��m�;�NZ B{f�IL�M5
�K+���_CP��GYM/���Y���5�A�p��9�2���,C˕];H����sa��V;+��č5y�T�R2D<��9����Rֈ۳G{l�in�?��YYY`�J�(P�S<¾��������PFgE������p紉3���;gu%o�F��B� ѡ3�<�ٴ�f��iPم��]�#]���뱈.N��7L��uR�����?QH�͑g��faW0>��$M5N�����P��AQ�`��+��ΰ���s� ��]�}
������>�fFs+̮3��]�p&navz����|r��h��.��\����

�i��BLNګ�z�Zgf	ܰ��è�mѬ��6��&���rs{J�h�kT�9`��<3F��Y3��2����!��V`�;�T����2x��L��Q���f���ڴ�чn�!RN��w(K���`ܞ�%.�,�e���]�Ȥ֟i關q�_6��@��_���X�2���N��;�+f�S~Ȳ�E����g��؜<��sǐ�8�� �Q���i�Ii��	���)�U�4��(����-Va�7�yG���W����ĎS���<��Z�����j.��m<ߥX��O���d���.z0���չ��[���^~6��z	���Gm�s���V����6
.���Vd�@y�,\���g� 2�t�$�12��J��o�O_�7�4��\η�f!�6!�����c�6�u��^�Lgy�I3+(�	��P����-�Q��L
>�96�1K뼱AöEw2��L�\���t��A`��8�T0��PK�I������:�_bđ>�`�O�Wq�=Bhi�C����;i֨�"Lp�@Fn�q�P:��Z�����Uܬv���bw1�<��[�4��pFRLp�qd�G�y��ж�*��zH�ٺIn̚y3Q���i�֛�<ՏZ����p瀕�|j�B���1�z���8.��:n�Ȣ]߂yUX��ñ������l�u�[��61�j)����;�ST=����	;���w##sϬ,n.�/!���D3S�Ӎ�v��������$�4	�
��+bNG��D����+Z��a&�#�?2�.j�9��
5K���fA)�m��մ��b����O^�a�̈Ƨ�)����Ւ���أ\�͊�ݠ���L�}V/����R�����46�]i����%�;z ��(o��a�&\�И���hљPJ&�w^*<ĸ}�BRKKK!�����$���֗^7XY�rN���wY����Bحu�7 �!�w٠�t�K��.-Q���H3B�N�Qc�[��AD�0|�� ��F"�z-��£YL�5eE�É:�y8!|}iڻ����L�s�z�c�:Z���eAg擟v�޷u�����O_�v�}M)������w(P�X� ����
�X!�J��Z,�]��~���f��2�d��=��wם���`snڹ	�;�t�M���|G�pN�T<��U&QLY�Qn�2�9[�_v ���upበtC.���*��u����Ȗ̯X�B6��������V��\<v(�?|0�ܖ�r?emr�:����1��AR��8��ܩ���OVPo�Qg��~29��2�\!�l��	Pe�"�hn��у�ќ{q��稡;i�,�[�Y������+�� ���O����6z����Ӷ6�{�nٿ��K�gu�ӂ�?Q'~�N��3�"3�m'���o�t��(�b�!������ܑh�����^��5�6"���E-u�E�,c����+���P��3�f�����m��W+�$���M9�ݭ2.��T 5��>-V���|;=P/�l���(TG�Q3
�nl���E�6�Im�&H�!~��{�Dl���&~����(Gh�5���i�i��Lz�����%)W��q�k�C{��1mITkwjz���Ժ���̧�D�m�FmT���!g�6sMC!�DD��>�-��Ww8!�leVG�fLX�o��D%���+�C�o��p�LBJj|�ZX�AY����us���o�����צ�Ǯ`����_}E�����CGr촹.ς	���<��i
�kU1���x���1�����95y��@��7UF���N7g3 *w���C-crlX�گ�2��n������j�+Wz������qf����8����a���$$s�I;0��;ȶ�Cm	�+>��[�{���`o`�C�J��G�=?�+fd�[�T/Х��sݘ��ZʣV�f�5�*`&������ԴC6���p�A��2�hE�)l��@���3ؘ�ׄ�Y�~�_�_����U����M�Zsek���&w���:�/��N���x�bf>�Oʹ��^�+���?d�]p��=γ���)��-�ǫY��=�5��gf�Xҗ��Jzo���b�t�~=����I��]_%��!d�� �{�i.dF�%��E:w��;=I	�8�ngh���_��D��:#�k���@n�ū��;W�Z��΋)��3�Zm��[.�3^p��۾י|��~�ɣ�hQ��u��8�h��><��&�r:��{ؘ����JL��_�R�9�蟇��Os�"ȈOk#"Z�"�����	Z�H��]�N��#ve�Է���j1�-�.��6V����>(g�.��#�׀�$�Yi\j.��:	��Ϲ�[y�Q4�[���*9�{�(�Z�B3S&���H��b`B]U H��t�mL���B��Xt�T��'��UҒ7\0�5Gzb_	�dud���ך#��6i��	jQ��=�?��������R זOOG�������������l�����c�@���v�+��U���,�m:i�y���q)�#A���1��hɞ�w�Z�z���f��~u	D�m=���N'h��-ى��a����h�����=�P/Y�z�-+�T;Wv��)�g��,��]��
�#S���6h:B��zKwK�9��YGc��|�;��:&���9������!M��{́޽ő��c{${r�3ߧY$ۓ��sV[P�K��Sݖf�W=��Ô���6{V���m���O�*U��Z[r���e��%�Lzyd���r"W���.$8F��q�ٟ����K�wY�ҙ.O���x ��)��V[�/�>��wF�S�?ASV�*<�,�6���ӝ�^�9�;M�Kľvf����H������Iݹj�o��[�~�5l���u������u��mݛb���_���kFIU<�r1b�a�<`��4�����|��j�<U�VB�J8Ҽ�3�dH�U��h1�4F�zӥ���0��B I��!�h��@��6�H5Ԙ����->�*���,]����h_�u:�bu��f��}Tx�oJZ�&J'�{���ӱ��������2y���?�N���ԋV׭���#�Fj�@U���]�+a��\V���0��IɌ��$�ѳ>��@��
Nz�Nׄ��MY]�3%�ߴ�i·hA�fFFK�,�Dd���K7do1��?B�@�Ԏ��}Tx�<����`����f˟�dq!!���!7���\�X��q����3-��m��hA�Z~B�IaR�fR"ҋ2/��T?��)+�b�|����k�>��T;r���lv�B��/���`�����gk��
>��lg<e�Cr��D�V��5��E=��H;��Æ�ME,�%Ӯ�K�@�rmC,S��M��T��U���L���S�N'��㭗��&H?ܸbF�.עqz����nd�t����X�]˭.v���H ��
`1[��t-X��,p�R����K��mc�����h�(�����qZ�������_�0�@����t���rt>�LNL�f���Y����"�i�=��8怴��
�������A�Ԏ|�m�˦}���_� �X�Z���Pf����֦zi�qL=��6�<Bf�	#H��߸?(�����3VC#��~����W�S�4c�_���r��"l7c� w� �)���B��6]��B�O4bzi �4�^V��;90�~^nkb���2R�~%��b��r)��I	ڌ�os�J���M���G��d�/�T��RR�b$���
���e'�爼~��(��)&@��H��"�R�t3E.(��$�-^�&�f�����b׸��9��S�����OE�;�7��������dP��G^Wb��;>>lP]�U'	A�q����߰*�3,o7�C�ۗ��26�$�%��k�9I���?�a�2v�)}������}�������땀N���bG�}�
���`�A9���.D0)[� ���~)�X�/�&Y�s ?�~��+�X����$�)";*�#���lW��7�`�y�:i��U^I9,�S��<�ɒ�p�/^�Xb��'��ns|]jO�0&�$ ��eۖݻ��4���D:��� ����u�u���B�؏����\��^��%#Sdb��Zo#0�G"��k0>�Ƿ�,w��0���s��c����fסdpc�/"����\9�6_T	E���q��3�gU(k����"ϮV���YJZ���2sT�C�|��[�����x���xց�� A�!�y�����9��LFԚ$Kp6.�ޡ$����*y�)R�znIێ��;��ib��v�~�9^t���{�Os3��D�*�$��)#�T`���sF$.�#Z�zW�H����8	=ذ�)�_ �K�?�n���l���\s��r�.c)H��Rﲧa���^��2ig���'��f�ң����e'�;P�їd����v�_���Wv��+���6
�S��&�Q������?�4:P�ΑIEl�	����>X��վ������=��Y�4A/��63����3�*9��C���\�� D �#8f$����
��޵w��\�ztG�)�e ���f�M�P<]*���:���8���m��̊�o��O����1�K��O�q-��i��#U��S����p!���_�Ut�/����̍�"h��!������}p��}�b�Z��'���d)��@��n<3
�~̟�3�ʲ�j}��Uo:�[6�����l��6�O����vB���H!�w�5��s�΃@���.��!t��ￃ<;0��l՝*Wt�S7u|�1�:l.�́axd#�ɢ�&�c�{��?����7�6`V��㚑�����o��8V��q6�W?`��eWd���P���꛺Q�Oħ�����q�0�� T�k�8��{xMk`�@3H������C��ͷ�}���
��-"����CJX����R��X��n����?��mo�b��8��#k+ip~~����}��K�a�QE�s>!�<A��*�_�F�{S��N�9�x��ÿ��s�4��rp/ԙ	ˎ����Zj+�i�Z�����ڒbJb��\&ݜ���X:��agG�E=ݗ���z��f<��~�I���mc~�"��������ZIh��%�w�zp�_�>t��K�����A��۪��T7���ʹ@�������cF�nݥ��d�^%�I�K�l^�|��D��d�U�BZ��:�|�[w�A���Y"�q�H�5Kr�����t2���c���pQ�2_��n�턘7#ݶruu(��v�ǉ����o_P����%��D���:n�8�p_2(k*��w\�I��_E��A' �矛D�:y����+b9��[�gLFG�U�4S���!�n��M���A�SY�����KǚO?���ki`���s���Xg�@C�������8��Up)E�ӵrhp�J9A�4�����_t��6�M+{'{����o���&Ã����6;�X���5��I
�c����ik/�ȓXdY��I����8���Cz����� ~�Ҽ�Q�N6��j(�D�~ن�4��Ґ7_O�/��{��ap��\-v�=4ۚ4��Z%�}�`Jw�����\�W�s~��S�frٌ=��Zn��q��.���6���b���QRn�?�p��>�0n�����bj�q~�
S��^1���l=��D`s�����&x7�%ν.�
���4y|N~!��4�� ��M��QeoQ�p~�{Alk���	�MX 1��v��`���H>�G������yԅA��zgpu�b!��b��22Ys�.q,LH	��@��QG�0E�Pt^�ӵ�k�=DN�,��T���恑���T�z7�~�}F"EP!.�O2��TƕHW7k����1-�c���~W�A��N]�;w<A3�	$�)�
 H����#�1��������bR���~33�4C7)��}[��_.. ,�D�^@� n������'�<�u�������߮^�$7U�Ys���ϐ��3�[���=�i6=������l�F��)BPWZ���~)�����?l��%�4�|�V�I o�9ߢV���b�
��i��3J5�^���KZy����HV@����-n��3��q�p�±����7g�CW�ޔ5J�Dg?�o�7ۤ�_����.(�����Oګ��K�a@F�+b�tI��L�z�G'��i#4�xkύ�E�R�ã�N5y]VG��J�N��S�_ ���a���7a�*΋3C��,J�ښR,�s�y�]@0��o��_�G��Tp�:���3����׾�&���[�wr�T�: ���-��S��_c�1�ҷ�o�<h����+�9�Q�r�PP�B�9���S&�ﻚ�&cr�-��O@K遬��j9O�=[?�j��	���q���3�eTgk�Ii�kl7��hg�q)~�y4�����i7�HS$4&_�C}�����F�w�*Vș9�e��{Z��V�������^g�%��i�&�Ǣ\��s�E����������%'�gsJ�5�/��z������5&aIQ1���>�5UP_݈Wj���o������r�	��t~������Ҽ���c^��b.�GU)�$�͛Sa�r7(�K�n[���'s�o�_�w�F�L�`������h���V%�!���y��?�I"�\,���{T��Rz9�V��o�-��q��t=��&��jm��k���&�H�<۷Mt�lA�q`����y���p����\�z���3����\������l���w�Ŕ{�RtmBV�ƾ���k�ə���:P�2�A�~J:j}_��d�;��������>�'�A �h�bss�q	�~�2k���2���]��3W[�n��<��z/���0�d1a���|h�]ck�o���y��-�K��`������&�J0�
�5!T#�)��9y��N��ɭC�dHs𻥩'�GL�Jc�����ip��cB�\(��#q#�mi��J!�qԻ�hW������U�0C��o�N�����y�o��O4�},ú>�d�Ȃ���z�yQ��L�<9��oK]>j9o"�rm����EJ�O�ޝ11����oe�����`u�OaBY��us���văl^�1a,
�<h��k���y|yDA~���%�ON��n:�ݵ+��mܨ��|fȃ�K�s���f�֘N�MY��%]$!W�?,BÜ���z+�feMm=��)z���?W�%<X߭�����%���gCC��;�wT�ؾl.0��P��k+<�l�PY����P� ��Z�G�7I�<�[�:�`�t���5c�}�4c?U������2���sD���㕪�[�QC}ݨ�3�G^R{��ͫ���r�֗�X?2���[�#8��M�뉞ku�k�wܑT�Ft�]��vmJ>~�J
v��^�<Y�IԄև�̪�H���ɟ��ƫt<6�����5ײe����3A0PW�F�Ҝ��2�^Dq)Tt����eI�X�(#g@<�m���QR11m[�N>�7�BJ��n�"E��T<m��c���S�Qb9`����O��LM�I��I�A���0�Q�����i�/��k{��2j������6X�Et)�kW|a�Ý�������{�ڔ2B����#���N�8Bv�n (�i�_�����Q2ޟgq��HB����պ��'dD��U���'c䃙�a�=��򺅘sª�2ƌ�M��h��Q�s�Q���-��:#���sE�����q��O%.�Y֧~l��1�0�#=���WD�{�v�::�m�>:*�sIm�&%�!��-�%��YN�!�t�����H�mWTeqr4[�K�Rq���WL�=x�VV�6	t4����n
��[l��Fv8z�Q�?���5�M_�=���%�Wr��҆k����#�l�(�Y	.�ӷ��1`!���b�H/��e�m��/%��֧>���L��E?�W�,ζ��7�BS]�4L8�Xtٚ�,,�T6�q>`�w�n�HB�����ș�/]��[��w=�-�~N��ri�#o��q�]�e���E>��(�<���^��c|��k��w!ۿ��;T��s:i���5i�l�/���ɺ��u,�xu-����<M�2�z�ɏ�%��Y��7�P%�>�ӑ��B[U��9�����`V�3s�$s�o���w#�$䣐�,�׻6��Y'\!� ϊO�-���y>��w�U���G�D��[]�_RK
�)�ӥf�f�FP�,�?���6��x,�܈ <��&4�E�k7��jx�.k�@�&��#����ՙ<&M-��w�cK�>�3Y����`w�6C>}�a����ugv�.`����P��w}�)�˃O�Bv�tͬ��������_�ɺ'����A�:��o�y��NeE���T݀�S5X��ƻ����iƾfu~�@�����<u������2IKK��_���{mB{�6��x���~��k�
�� ��5�.<r;=��&��:Y��9��I�x����CnR+E�m�61���������%��\�v�������U1s� P���8U�[��q������~/�������Njdo�g��8<��SB�r���{��@[���� ����?���j�X�i��z�kt�_������
���teC�#[�7S���1��O�|�S&x1jm�c�yZ������Q��B�3 G�OA;�����X�$�hJ����T� �z�V&��9���Q8&��1�:P�p���Z�<v��t>�7��]ko�'�RjBi�u<�E����l���
٦B�Ts
���^=�=jM��v�����;zbd+�lJ]����s~�I��~.V�k��+�Ԛ�l7�\3����.c�<�9���0x���qŜ�����x:/�r+���%y�.���ￕ&�R�ؒrr��,,�QѨںڒZ|���U���c<�ؚ���З8�^�e�[��p�Ѷ���5fE�e�����卜N!3�t!vQ�`pW �֏����S�,��Ʌ%������h�KK�_h�R1�ejVo�<O���t߹\/yX�M���loE[�s����R:�n2�5����
�Ey*�.3=��y��Yjj��diT�[��"pQ��3���6�z��T^�RG�E&��d��N�V���j�è�Jo���bs� 1�7~��7�ـ�69N2��n}�ʠP�H$/�ī���ɽ�h9<P��n|���ooK�V���	Yuݹ�V�o��LE� e0n�7�18�k�*Gp�t��PA>?\y���m�9�Fl㑗�C)���q��"2t��Xb���i�=|ﶶə�P��#I�I*81������N�����}��F29�t�W �bb6�vr�>o��> /�j����!݇���]�].�HBw?{�.�^����0�?�9������Zym\�ڳ�0A��+�hȠk�����j���M<�[l�i� �G�<ې� ��_	���xT5��H�X������0؅)��}I%�yGKK��T���/�R��,)f��1�e�r|f���L�IC.~I�$k��O�����rG�����$D-���B�h(�Dml������R�=X�eqab=���[z���n���}��pX�+~��x��������j'/D�q��R��7f��M��)���G��f�g�s�ޅ���=۷}��G�	}_~��`��BZ����t��,?v�ɷ1`BR�.Nsg�˘r� )����~����3}��_տ�vj�E��Vw�и�^�z��FI��:�0zO�,�z"u���hn$�ĿQ ��cQ�+a[[������}�[J����H������р�c���{�ِy�3�����L����`٢���I��)�ZѶ-z��o����^����ң��·
��Dc�e�TD��j�Q-��H-�؏��j����Qo@u���'W��D�k��Pj�R԰�������a����(�C��Ad��w���j��xQH�U��RDj��*@�\J�tn�}2fD���WXI���+�>^K8��9Ҙ�5̫bb�@dK�%���A��I{��!�h��8��ډd|�dۉ�%����$H�nԵ6Y���m:k�:r������ى`��s~�Dy�W*2�Y��U?"C�B����+m!Q��nnn���b�w�e��Eߛ��[���ܽ���	D|9=$6���~�������+OG{3a6�9 �ؿ�s���<�:���1yvs۠�䁈a1�4�����a0Tb+�D��	·� ģ���}U�#����éA���r؄�O´Ԥ\]y^:�v��r�py_k3IK&��E���:V"߁f:�%���z�LD�Uj&M���6�>���f�k��nsU�Ƭ��Y�� y�@�#������%֣*��6�vB�����N�֚�+��������9��� �F�-P�� �@O�0��ӓ��Cqa��H�A�ȄM�]�E�RO��[>��k�R���f�Z5<��p��B4T��IH<`Pe��{G �vDX�jwEA~��{�ܑ�J_u�;���0X2�>��X��D(^A^(�ݩ��闫FF���Y�M��x��?�~��	łY�kD"���y钥Jl��\���)B
LG2��)��'0^��j�x�G8P��Ҧ}28v����1�{A����IFJ�T���@BBZ۹�^���4���� ���p"ŵ� -��T����!����~�>|47UI,�m	�C����|���$� G�m���>��;��XF��S*�������&�У��� ������]���!�?����EoVC<w�<Z��5���ns/��г�����*+��{TM���K�+�z&�����'h�l���:����&���_u�1;���2����Q�}2�@C5@瞴���k쨨���),�C��:�~qqaz2��;��� ԙ546Z�}%��m����mhj2�.Q�m��5���@��c�0R�+$�W�� 2ۏ��oн ���`�\��|9�BOW�t�m�ԭ�EG|�jʔ
�X�M+�� ����f���^�ڬ�e��W���L�+��XR��zH�h�=�'5c�{9�����A��[���E{
9�"8�a�/���.�̨�*�؏f���H��,,���=:)�:��KR�̩+��]7�SVs�5ɬ�����W���;�Oe�#M���W�-��k���BLPo9��{Y'Xq��8K�;�-��pZ[O��8�^�����-�|����	ψ���H�~�ֿ�ϙ_���!�r�{�6 eˁ�0`�I�к!������թl�h��������3�5���+�����s�������Q7Sm/U}y��t�Q��UPh��[b}�u�����w[e✝wTj�"��Gߢ--K�9^K�V{O{�C�>/C%���v&A��.�R�$ta�a.��Xr���
j�Z"����(�j�������k���i��֥*Z[[[/G��X��CD	�~u(��s},��*a͚��G$L�7��Ԃ[�l>;g(`��bw����֔����y,r`����1���\����y���<�ix��M����+��nŮ��d����Y��+����ى!�h>�Ǽ.���@�]��g|NN�K��"�UTa�6�AhE��
#�hDe #K��}G�t5d�}���R��[�Q݁����G�1c(a$l�9�ts1/�����l�[��||w^�'����p���p((�]��,x, �99�hk"}�U'@����t��&(�E���ϖ��88��uk2.Կ��:,baa��:���� R]����"�����Q���n:� �t"ZՉt�'C2ЇP��ֶ�8�G!��R��lmp[O��� ������o݃i�A��:{�6��cҤ������P���nӐ|۽��Rot; �*�@I��Ҥ��!ߓ�j4�o5vKQYd�M��,W��ӓD]E�7���}�-�����#b.��g�4�).�M��:�FB�D���±�Q������6��ѳ`q�QPJ'�~~J�{�=��3�b"�=nLs���<8.i)�DO�9� ݎ
er�]>��[�,�B��#��o�[.w��;�����$�ߟ�f��E5�a�G�-�m���)��~����}?�|IWz$j={�_VZ��Z9����N��5o>���@��]&��6q�%$�;��vt�uIc���d��0��cg�x�#�|����mh���z�bd�Uo�F&����,�LČ�P�`k5���SmG���ҟ՝Phjz:��d�/���0����t$�����KY{049��_aޒ�'�'�xOw4��Ki������`����r iU�&�+G1W����U����� �+�e�܋���cQ	��Hb���.wG8�?�­5D.[�b�B���s��Ė�Ի����W�W��@퀖zk��N٠�o_(��g�(��g�{�3��A�6,��8V�8DA�\
��G���]<�]����	�p�\A�f��~������^����;��@��Zw@,Byhd����nt]	�IrugN��tS`C�x��gY��2,cbz�u�����ܳ�yKI�:x8�vg��V���'79�B(6�XI^upu�Ĩ Гk���>X`Bp��C�2�Á���K��5�����D]2�RM��u�J��<�1�f�aw�� �S���kg�'`_�nu&��e)�/�U���GH�iao�!-�&��_��)���h�q#��BgCl�	��
��@r<zy���Ef{L����ME�Ҹq�K�,�䞣w��]F^E�(�U�b�𤋮���Í`��`�����|��������&Я��0c��2��3����}*n���K���[��x��WРұ_4O@#��ӊz��S^�5 P�j��CD3=�;Cz���*�xߪVM4P���np�Bq��O�u��)/�)OT�f|�@�R���-Jv=�v#d�pW�� � %?/�VA�u�.����&�$�`��#D3�P��t��㊄��B�1�����́�K����y����/AaYș8;�<��[C���{|�uύ���x����l��r./��H.2�$M^���}�Ŝj��ٶ}�IYv�E:k7ϳ?⒱�)�id�~�������/���lm��`
z������q�} ��8���u�Y�o,}"4AU��*��Yn��,6��^ɩY"�^D�3�Q7W߄.���9.J��Fs6~��:j����UV���V���[+��ot��m:�W��M��<�E띉�b/�I�S;#�J�� ��\�B�<'�A�ir��Na�����煉l�K���ިפ`Ѓ�U%BvE���`,�8n�W��#
߻�RO��)��H���y���ђ]Z�t����n-��w��)2��W?��A��'����^�Df�����vh���P��K��λf`wЉ0ܵ�
�=Rts��2a�r�g6�ϓ5AB���6��N�	b��B����r�n����/7NMvH�@&}�lL_���(�
�v�-��2���L���]5̿bDV�]�_Q��с^Ŗ%X�	91J,I����Ә��_Ϳ,�X��*�![P鉒�t<���gy���|��Y�s���(a2jh���9( ������M]4A��B��s GuǗe$�~��ٟ����#�.��c�$Q�O��"��:e��ۍ��;�M'���+�+�wگ�yZ���&�|��X8�_䉼~��ް�v��xTn�3�[9hq6�̇��r���� '��X��I�L���W�!�SDJ?ck�	mS��\�r�[�z���(���eu����AFLr���k���[X=�q�0ø�c��H^�v3=^��<hĘ"*A����Y��_4��%y�)���L�*�q�m��}�n�+\�F�����Յ�|Y�k�(��n"�Q�Au'E�)�$ "w[W%�8u�����Xf������LIG�WM�/�#'Q�ۊ��)D�� ��\|�7�T�߬����r���L��>�,y�m�Bs���Z�L>k~l���oL݆�6�@�9�~���Bd�gu�q�l�c:���3�j�m�c�ms�QLKo�����'��&鹫��O��"�u��W7�ޒ
�3!��U����`P����$(�ԉx�򡨵
�mvN��:��͸;��~�~��@��W`���t��W
��.���E� �
&��G�������:���vG��u�U��P!Q�ޤ1M)!(��@���Ӱi�>Z����D|�_�Uݵ1�2���і5�&����]�}�+>�.ح9���:��N+�Ԍ����x����p���ʐE�7������P|�8;�\�=���0����	���Y�������3P��VÞN�k�N��K���F�W!zЈ��:8`U>^����|��9913�e���~t��%���R��J�|�] �u�P��ر{�������� �����C�in}mG��������y���/R�2�_��>},+���Q_�#������N���j���h�[LbI;����݃2�u�4Jo�nsʜϭ���ytk��q��g����7p�xU�,k�%'����R�%(^nJKy�	4�1}Y|HZ)WM����n����@.]Q�"2��Դ����=:�LI
�����^!z�~R�̟"V|���U�.grwv��8,X����?����ִN���[���$ʒ�H�yR׽�`53�����5�p�ӓ|7�s��z�m�����i��p�`�g�U�|Q��0�8�@�c'�F�o5����pWӑ?'��]hO�Tg�����1Ϯ?���0��޴~7�h|q[s����m'�p9�l|������k6fV�3����h�A�T�&)���`�	��f�ۣ��$�IcL����:0ȷ[e�Ź����0A� l٘;W���n� F���]Ȋ+�����<��v��Xw�R�J��SB��	R�s@K�]��'�~�T�H���]�Ϣv�d-C�.��j����j��k���}�_��Ү`G� dac!:��XTB�?�ţ�Uh3��9N�5D��=&��/������-}<�5�Zc<��9�*)a�v�_gQ�쁩�ǁ�#���icJ����$�"o~�����~=��̡����!<`cv`�z��?��"�X_U61^:��w/5�:��y��֊���tл�z��朊#oo�ɖ��86�\��0���V��C�wF޵С�D������yk52���:�����*��1	bB�S"h����zI�P[iO�����E�D���/(a���w��Ƭ�g��tl�Ӎ����Y���ϑzH:W��6T\}	"�Y_PR�����)�g{����AtA���U[W׼?ՖHScW������xU�.�	�<o���
I�ֈ��**��t�~-��8ώ�
���� ��Wf�c��n�4=��"���*XF�u����[�$����~��\j��!j���TLd���(��R2���΂�~��ɉX	�t1[_'�^(�P�M�Dރn�)܁�{�Cz���`�$Cm-��TW\�8�z�16��!�Ђ��Qv앸��"�W��,nn˝�A	��OClՌ6���XȺ�=4�q��x�i��ZΈ���:-���(H|}�*K��l�a؄��1�((�-e�~�7���%�	�:����@�Tc���8h�7���E�lXz�
���r�Y�8f��+1��n�O�$2D��~� �|�/��p��K�CJ21_�1����rs��^q
��Pj;����j`�_��닉�E�G�i%
hd�uƐ�	��H��蹜����-���Ⱦ���Ͻ�jW/�}��oNܙ3�N�7�ĥ�$o�,o>\>E2���[�Aq�0$3��Ǒ��1WZt�I̋�3K��|�>6]>��=���Cw��&^���ZT��?�H��Y"����S����]�7Jns�+��C�-�6A�'��FF��%�f�ݏÐ��P����W;T%���B4�:���Eo�'�_�?�.还��~����r�1(���ɻ?='�����dm�;���U�lY[�����m�?	1��G6~��*z��o�[�}���pq376��1Ŗ�ª����"��!M
X�E~D���Z�e)�y//j��/ו�i�U��ݲ�jH�Ռn����P8��M��ʪ����'�כ1��*1���A��=�4ڦ2���j�F�}02�7_g���u�����ii>(�rO���0�)ҽ����9�&k�fub�ڠ�8H���ᜅ�,���Аt���5����A�JNx4�J����)��r���Y1]���va���Fp��A�<	))ࠪy�A�6JG����w� ����rl�MlUVxx|�)]_p�?�U���!}���W�]~R���@�7a>�T;_zQ�Y�2��.�?�_��������Ø��z�&q/p��M�Z�h���tTP&0`�q�n�9�.|���� �:P�$�N9n:>���`v��0�W��B��Q�[Z�y�
k��y!Wf}u���8�馉s�
� } 1��ݽ=)y�c���"����EL�Z|�,XP.7~�Gy�q�gu9s���u���7#����H�-^�O�������s8�o��$��!f5��qyh,��a���W0�+��M��R���I���K���T��ddrKKb6���CE"i-�]B�0�4�B�/4�{,�E�P(��O�X�Y���Gya�	�U�nK�c��ۇ���,���I��ek��Զ���+�E�'�$$�G�����|��8���7�W���9�,�hi�䷥qh�HnӪWgs�>6,�ik��[d�,�cHNC�rG��z4�DTa���OX�S_(
j+��"=<]UD3K6��{�ַ�?ؘ���Uڃ<$b�2|�-"�6;��,�KW}#��C$�Ϋ[�0F���q��P���-'�{�)�NA�yE&ވ�V�b
��)���6��R�6t�<Utii�����Z�t�!�O��{��ق�����&c"����Z.t_8������aV7�GS�(��,fTo@<�l�Qz���K�����:�f�S�ӛ��jE����հ��1�㎈
�|� {�m2��,Q��4�H�0���xi��+�f��1cϣ,�GU�uڼ��� -�F�;<�I���7���v��Q�/�Tک堫٦î��#�q� CA,1�~�B����%�a�>����؍ ����'yT�[A��"p=���ewW�r+�I�6TR�
)Z'+���b�����K��q�8�
K,8�t�V�A>�wz:J��	�82�r��q��m_#hҙOA�����;��k�d��F�[8���
��޶����>)x� 3�]��ǿ���>�>�S	v������LN�П9�aV�	����:�̃`�%FW����4AGG����aO6��r�	$aџ��}۷h��NR:˵Qk+T������ފ�u����c�T�Z��Qt�0ij�l�w2vv�e�WėY¹�)��H������i� �3s����Hc��f9>�#
���A��/�L2�C���q,L�);�c̉����@GC;�E�����j,�����M7eU������6��}�m>�z�r ٛ��[�E1�a&<�?��:*�����S:��S�.I��隡�SD�AA��ia�!��!���{���5���ଳ�����s,���·�ArA�7A�?ҏ��k��F�X��T����'d�Þ��n����]]</SLL��Ŭ�$��o�&����i���[Wv�"�Q�d=K�
 ���/݂�1�ۼ:|[ǥ��W�v2u����u9Y��u���w=�vࡪ�W?^EU���'Yk-��\]��sw�Z�x�|�@�����;{Z':R��~?$?�JKKN����P�@u�޼+���k7b���#�h���OMV��g���}�viݧQ���@1Gl�0���-��ڮ���L�&;	_��p�nl?Y��-�]��/Fŗ�������s��OKio�U�;��Z}8�k�gn�ך~���DZ�h���j��*EHb

�u4I�c�&��׳�lmK]��gA|�+��BGG�ւ=r�9�GE������3;4E�f�ŕ��ۿ����1�ϑ��$����������_
!��&���Fh�Pq�R)�l0���Z�u�⽞pu��x 	UaN�ñ�WN�$rZN�:V��y �p�!�ig!�0���G��*���Δ�јe�ϞKp�͇/I�d�c;��	bEU��R{�C�kB5�Zx�Z:��ӌ��v�������-��.�V�B����"�u��9>a�zZl��{:�-��F��Ġ==���.������]�YI�?�����Djk�>'�@/��ʂ	v��/�����X��U
���;��I�0Zt6�}��w-�dq0���m���/�ϛ}ha�4sE�Eg���V_.$�4٦��_��*1[�=�o�Q��>���c��P.W����yj�2�NVv���b���Y�W�/"E<���L��&4p�w���|�L�Th=��!��C<�@ ?��4I)�i�r@�Ԋm�}��{��� ��f1 �d�$D�~����H�?&���,�$����Í�d4ùJ� #��-��E�?JNK�Wd�s�G!��ݫY�[ſ�Ԛ�����fP�LS�D|�}M/r*�Z�uw���v��X�ť�njW�Ly�Z̨����¸���紲4�ӑ�"�vg��|��e���L���Svb�߆W���WP��oT+��0rj�*kj��!����[�����A0�i��N�Z����;�^[��Gi�N��&雗�~�T�ߧ$�>\cz~l�lזy5_��w���	w��9��.S�x�$4�~E�Qa
�r>��h�4��܅�K�*^b��d�?8��Tֶ����d>���8�&��3�>��2W��vvj�Xp�!>ٌ-�oO���'���a%���10��AW��$ؓ[ �,����%��J7[t���c�YAi��f
+(�*��xr���6&C'�)nw�}^�������k�$��_2$�=�%U�������1�;�1h��˪G�O!fy�-Tn?�c�&�&��c����6��r��)_�hSK�s����Aw�䃣_�xS���x�˵B��k6�3wyRHn�^��p����^�����u�'��5�K3����+��;k:S�;?nV�X�fB�����S��90�Ԓw�@17�t���^�fg�{D�n40'����WVjv�BFh(:#���$�A�:��ظpwC'2cu��̚沉����&q>�`�JAj¤��F
������ �9�	n�$v��g"m��=+ޏm�+s�������+��OE�W�j��0g�WQz,*��b�ϕN��
�ʰI�
w���G����gffĭ�h��^�9%#��)���J�=�f�N��6C��d���?�����E�;̐+�� ���4�8	��3�C8Ҳ;����F|���3[(ޟ\������g������c��^���.����\�=��[�rov���(�����Au)��6�d�Z��N)� 7MCl��� S0%�Ve,���:�Y��sa��3��L���{&��ߌ��{v 1q��ʼ�fܴ�]A��4>ԉB��r������	�	��Α��>�k�6��f�&���^��:���V�_��Yd���h�v��N�~�6�da+�j��.o�����E��+v���k��Si�8�r�К�P#�������r���+�Y�g_���[���Q;ntJ�g�)?�gǵ�Y�.v��c}�C|��ɕ /Z$�Ci��lz@A!c�����{՞ns�r%T1��״��pW36��<�g\IҼ3u���t̃�t�����L]ڰQ2�ݘe!v�\s`k)���(9l�Z6Y��(?ں����iZ�����Z�7�Gd�}�ж���JM{�y�'�D���"��=�\��f�`[k����{��W�Y�<U�D�~�������z6,����n3��� A�[؅<7�+�ܕ��=[�
��<�ʥ���y�*���i�Eȗ�zng���g�#l�pz�2�1:Q�$aX'Κp�k���=±�΢ҍj���U�P�� +?,w�!�ɋZ_�����N�����	�.���n�W����4�����2���>��\����=Wx��FQѹ��hv� �<�6+I�a'U���,��g�sav"���{F\��b?�*��{����[�GY�e��pw�����1���n��N�տj�-jƂ�:���-1�1E�G	�ÁQ���e����ʆ�w/�-��0�q���V���:wa��g�|����y����-̰r���t���`؅FXy�3�����sЧ��[�;��X��Hk\�c��>�<=ۭ-uA�1�I�J�x5�a!U���՛{^�Y�e�3I=�w*��.��i�?λ�Af/QY�7�%3~���yv5I�[W\G�$s����4�~�RWUH��0�
WCZ����G�������̆[Ƨ���	�[i�-n�GxD�n�*��<u�H�5�\�;�\	�{�z�O-6Em��j8��i��ꍍ��7Ű���͐�����E".�Ń�:TdCqdy�����9�2,����'_uǿ�TT�H.����_�+����}��Ӭ��_B�յ��4"Ʋ���"gB],1���x�'����)� ��u���)͹�Dϓ�5Ӭ\]�KO����%�YM[�3�	��)G��:J���p��L:��%�c���Q5"�9w<�R7A����xn٢����"��+Ո���5f���@�8B(b�2���p����6�o4���\���@̪��/���<����f���w&����a+}�h�ڔ�m_r�I��t�%��3hG�d�Z��u�p�˩�2��#��ۻK K�>�qK;�D��&�i#$�E����V߭�'��*��*�"-���h��t�A$�pC>eU����p��Ap*�{)����2W���*q���3ޟF7[?�O	�C]\j��t=��6����ͫ�����X^k*Ə���,��\'c���B��M|��ZJ���`as���'\�nwvb�F��/<e��A:��cU@�2��=/�g�x��~2��8�ֱ:a}J8��g�$��)�����m��,V
��2}�'���b��@=��om}Z��έF��F156�[-'�������}2h\��?١�O�00���g7���!�5����u��b��)�+�$C��c������ȓ�� �ZD�
�#�g����Fr/��u���(T�:����s�p�[����ëa,����E�q�7�$0j�p��H����
�Ȼ��OZ/�v�*W�^��5�[�B���	�6���"z��cR�1��XB������j��l�<�� k�/l|�t#��W�͎�,nV�y*�
4�Xlۢ�$��U�m��}MC����_\Ot��������>��g�`���b����_ʋ�\�ܸ�ǯ?��Hx�Ny?dڞ��Wu�|�Pc%��F��;f��.E��ty'�Ɔ����|D�M:�㔗�_�e����$�I��+���,���̾s�p���e�k�$:|LT�C�K�)��������o��.�| �flՄ�29o7��Il�����s�Ћ�d���zM��R���?k9�'ö͘�$����M�5i����[�����'�?�@}��m�w���K�lbkŹ�w�l.�'�A�W�?�S���>�?�2���0^<���%E:O�뭁'�Q\%�%��j���x"�R{�a��w)��l�.�3=ny_��H��	\�Sz�����7��Ч˳��\���,��Tm��f,���V��M2g�p2[�'�������
�N���Ob�/��C�/����k�3����>xŖ�3���(����e�����6�3{4J�/��h�iDy_��ʈ���W5��9�X���D��7��2_��h��@;�hh�9�*	`E��@�X�|�H֣��+M���1n0��͹�H�|�E(1���v�����n~��D�m��Ʊ�4�;�y�>Kt1N�n����=+��Ý�e%Ohбw�vk�Ѐ7�b�b�(�򂶵RYScH�Ϯ��	Q�p��#�zV|ZVܼ�;Z�`�+*�F�ɩ|�%Xd��;L�����ӵ(�! �vM}X���\��X��yJ�����u8���6-_��x��s���4�D����[��1'����hc��%�ធ���&�3d�sx�1�W̧�) Q~F�V���m�7����ϕ�_�d���_���z3N����v����q�s�-�V���d���g�+jڋ"ĕ���=h%� ��B�A����G��������HG��v�5yq�-7���B��r���9�I����)j�l&����	ξ�P/���C΁�sXP��ŖI��E��9��2�%'��`v7H_V�{ǅ�w�L�*�Ɣ�>�t�<K��g�uq��*nr8"}�~�{+\es12��T�I�8�����8���qI�Ut��#+�5�y�wv��k��0�O.�n���V��l�//.e�r�������r�$�Ɨ{�!��h��.{�G���r��?�]ޣ��9[�Ns�[�_����);�:,��j�4��T��~twy��ΐ?�a�r�t|t*��{<ud ���t���]�n����E Ua�_1	�C)ف�b��]�Y���n��XMw{��å��\��J�~����$S��eEf���9�S�ɗ�M���/�>�I^)#gI���=)p�]DRyV���sW�ĩ�q�IasZ���u.�Z��a��X���Ј���c|�b�O��K7*性��e�Ҿ,k�0䚥�|A�Ҙˍ�}�KU�t��m���C�KЭ)I�'�5W�}�s���9 ���=���[!`�7fA	����*�`l2��T-~<F�_Fh0���%#)�Ά�Å16v��w�������D�Ify�C~�1�JxR��I$T��	���<3zv�G��������ox,��{pPna����5p�υ���ur���AXK^ل4V8@��79�B�X�&^���_PV�ۥ�9;��&�Kc�'������S��Y��\����jc�*I0+3V��g�j��K�g��]8!B�E�	p�7�m��<Ί~zlɾ�5-�d	����O�YvM�>�f����靆�Ew��[ޭvܲ�-WbouZޕ�q���%� nWҬѽWW�������,I��w�Kw 9��=��[��2'�xbdϑ�������* ��� ����������U�c��IeKO�|BN <�4���q����L\��T����2�~����^8�q�.RV[�<���]`!E=� �N�_�$�[���,������	<���ht/`'���e������R[�1�-��o�"*�N�k��+���ٓp�D��M��ɕ�#�g����vY�VW�D�����Y���M�B�$��W����>w�a�(���T/@`���B�84gزeTΑ�K-��.ǃ=
��c�pT���vt\1���5�g]�������G\�� �}7(7���̅	�n���"�9��/��ik�/&!`Ӻ,���,v�����8ƍ�q�>C�'��Z��P�����J	�zG�?ˁ"�Ν�#��9-�-��R+�a.G�}3��2u8��9�b�_	[�p�8�H��-�[�C^���nX3+��9Q�O�o1G=w�J��[�F i����~���PB����8��F5�V~�:�b�t��Y���e��*+������Љ�Y���=^����`V�O	��+��X���
+�]$l�d�������� �� ���Ȝw;�pI�u�7U7�Hw��{�?�Q�ʬ[���/ex�����q�� W�vؽ��&<z�o���ۚv�[=�K]�]�@���Eӽ�_^�<��>T<w\b�@6HÍ/�I�V�F���KGW��6~�����hi�*	\��u���uM���Ž�;��4_�Km�XMz|�)[�[nN{���O���i+�/z^"a��~d��L���#ٺ�iC�}o�<�-�W�N��;8�}U�ÅS�����7�3(1�z#� -�����p$W��.�����H�AK��Mn�`��bO�4�1��ٿ�5������d������p�4s���Ɖ5��c��X{�Fi�cc{�:�B�{�fc���[ �p�,ꅘ�G��L�W��	~k7��|ςڿ�5~��~i��D��������Q��2q���mA�Y�Wl���ӳ]}���(�)���z���_W�p�IbJ���U���U�}q�U0/�n �K��O�/�e������zl6�n`	N �iE�03�@r.�Pd�+�b��í������e�5}�ajby��z��!�t|u�	0�+\�ѧ�~u��eV��i�3��ox��(=��V�o��Vצv�f�㯱Ʊ1���6qS���k�h�� �+\nmq�r3���/�d`������[���ڱ���B$���~��k�Bx��
Z��źZu�W3�r���σ�m?��Pj�=[;۝nv]{>[e����f;I��V��4b2g�U�`M���&�ľ[Dk�����d$�M-������A �\�����ѷe��证j$���^��gU�&� !�&���Dk�@��}D��ٞ�UبF��!�Ƨ����m��	�sL[��H��I��W��Y�����*EA�X*5�a��{��u�;aϋ3�|ˮ�&|��r��HD
�k�fp1M����4�,W泛��&)�Z��;nEn�,�­����	̺�I�6&S��	�gA�D+5������rL�mv��5�|Y�_{\��A�s���^�gG��h��}P�]�W8���Ջ�5�*��-��'���.��Z���s �S����Stt7�;A$#��&�u�G���[��}HT���(�!L�e/Z����H�_��{���%ԇ5N���W�IyI��)Z���O��J�b��>��������R�K������\Hn���z���G�}E�ihf	��	ש��="�p�Bu��B��]�pX]�y8v�/�A�@����X'�M^:Z�r��*f�T5�@f4��!�y����d(�LĢ`��a�k��b�+��%�+Q\DfT�e>.{?͂�
0ک��J���x����8�ؚ��3*cć[c��?�A*)�����a�������6���y�A����zE<i��U70!��I���!4�Hw��4��ݣ�;���;AGN�ֶ��M�ogg���X%955����g�(�x���0��q��冱8X�z��f��{r�>_��Ķ�1��y�m�`a�9��lH�8D[ϓ/mh{>�$�����ً���Lq^��ǒ�t��:��.�3�d�Ę?�K�YU����ԄҮ��'K�'�����-�5�D�}
�t�pC�'M�0@�"ڟ�U@\$~EĬυ��&W�b�����Zwor�_����a.{,�z���zmXJ��,��x�˂��cr{,�()��I����}��'���[
r�OCK?Re�~���w�N��-s�X�&�8z�h�~Gơt}x?�v�wYg=�z�u�"2���%;}D��l���~2[Re�`߷�RjWjk�8�FiP�+N��5i8P���]]t<%��z�&�3�P�]�4����׋=H�֘�hW�E�c�p�/��ċ��˼��%�+;��Rlۢ��CD6�T4�2XE��o����t'��bg�h�Xl����<��J:���o�S�CI�όJ�+=V�.���Bw�b�I,O�gr���,끫ID`۟��@)�걟͹��1�[��k�u�ہq��|u��|���A�A��W�L��T<��ٟY$�B�7�ᔔwDVzuYxqx�A���dalln ���d	�'����^�-j���޺ݤL��{Pb@n\��6�Q��+e*TI�Ӓ�H/�_)����Z��p�O�����?����܈�V���b7ĵtcW�Y��6�9�Oh�2=h�u�F�a,���I�K�cZ�c5����s�I����XD�5�bHٟK���	Q�b��PA�%lXY�tg��c�S~}� ES ���#Wd	S�if�ķ����gY��I��\�
}2S�R,������P"���F�(3����m=���"���ʋ����Vg�~�{�����j��ô��?����h�"%�������Ę#TqK3�K�C��B���q�so����p����v��,��Ĭ����?+hBK����>�Y(=V��MB0��g[��r�Z�P���8�L{��|�+�'��;�98���ߣ]�3 :,��7����2��*�ڍT�	F$.J��mJ5���gJ��zpaU�zs՜��\� w��M�֥���Y���kL%]Ms�?{/t�7�Z4�K%)/��,!��|B��~�y��p�)�F+%�6z�r$��y�X�ȫ�osd��"�l���7f�V+N<&����q�q>!������*��8���1-`Kx��y�&�{�)|�g�J��-Ye�[Q�L��;K��.=�����G��$�3������
�hV��n��-������+ss��-m�o�a4����v&F<ݘ��vۍ�ia{�U)��g�	,�>D��f�
e��gPdVSp6��_���K�� �����Jf���7��� ��6N:�Pe{j�
�/�B�>��p���~�KZw4''��R%����\)�W4'~���Z�.�}���E@�_����a�=��A�k�>c[�4-n��S�؋X���{�x���a��4��"�7g8
�L��ؐ M��B[��VB��#�^��b�5�s7\�U�c��B5gDh�\2l�V��<�U�p��7��� _����*����-�m�Fs31R��5?�:`_��.Г6!#�@������u��P��xNω��$�ʸ(�E
��г���eɓ!C�"q��z�V��q���A�F�����	����?��ݒZrx3fV�s� ����5R y�@�������x,�&����Q����	5���#�~�9Ot��2��_��ܘ&��_�YG���"}�'�k������_� ���19oOv��YX4/�98
�B��g���b5fϾ���:~��9r �qB����'1�]H��b�����XLL.�9.Ķ��g:z�����L��R�}������7��4~�h�Qi���[:+�#;l
�|��q�������2}���W�c*�~Fd��5X����N�#�B,��W���~��/�����P�.��<׊�a��;XeM��6��� ���XlW0 Ӫ6��U :5����gV#h4G�!R���lc$`aʾ ���ί�u?���K%Y'$���>S �	נ䳺`ᣞڎ�`-�w;�A��v ����F@H��f?='��׆�^�sꏕF ��p�e��N��]����lWИ6Yʤ��
�@<*��ῐ���޵O:�~WR!i�1Uv��WG������ŉ�z$�n����Bj����o����!����ڔ?\�ߴ�] c�2��O�P_䌏{����ϟ]��0���W�7�����I���څ*����!�!c]���7zhl�j���	��R�A*��~m���^*�a�+��>�ja(���X��NX>�N�xb��aA�`t�.bsz�:�"����^{��;vZM_1�Ç�$�vL�� )!�yc5}��W:��c�JM�k�����VV���27�t��,[I l�sr���q3�Ek�f\���Y�?�@"�2�T$�Hbig��=���.�L9�}@-LLe�DZ��^�#��O������Ո�w��v��2� �~�:B�-3�^���!�ԕ-���`3��C�N��"tAg�A�EVY�B��ҝy2~���\�K��㱗,�0{�}���iʻ���;���2b1���G�ҿ�ʹ�8�?H�r�GM��g���	�lP�  ��/�/z��2e�^��3�$gj�K�8-�N��2.����ђ�! �(��y��&ǞN�{��7�ק>���ݍњ��[�æ]|�_�tA�����A#]Ɛ[*w=,:^~H�G�A�gr����a*�űG�mZ�g~\��^��\�H,��4~e�w���rqȺ�Ե�ޱ��R�F�`��ɦ��-`�㭅����3�t��|��}B-t���G�I7p��
Vm9V��iaI��?� ͋���g��_5�����cn�1u?�����ňk��E���q���;@�e<S�_��O�Hh�U�ڔy:m�@/V�ߖ]�O����RD탣n$�J�Ԉ�u�J�YW	���=��6��Q��̈���e���\��=P��[c19���*��z҂� �:�m�ҧ�v, ���*�2�q]@:�va�F�K
��E|V��~-��F��i�ࡪ�x0R��ߊD�Ws�`�F�'T��|���������9�r��_�T�~����q,Q,r9G�����w��I>�G6���K�wGD2X].��ĳY����Xۜ���f�z��K��������!(?|S��x����oTR�"��~�,�߆�Y�{_�l��07��CQ֜�ќ3v[n8⫆d)W��1�m~n��;�������X�]@��8���m�{���x
!�|Z7zHsQe����o�14勃T�����F+Xح�v��>����Ԥ�"���c�i\�-�����y���ZIM�
�������_�UEG��	���Dڥc����3W��F Q�)nS�G�/���e"��m�tj�c`ﾮ-�~��%1�m
��o���r25�'y��9�~�S��\�$�KE� Rlc|��{S�Ŏ1�lًjĤ��X�ъ���N���1�]J8C����G)�=����ym���Q�0+��lϧ�+����9�Ɂ"Z=Y��8QpLR%����p����6�|��s��Y�������kr��L�Lrr+G߰��߽CB�2�W�/����_?����o����^�I0L)Zcuw�X|�?U����x�0j!-ꤐ��BOc����\~8��h)����~�_��&h;�b2�F^">�^&�,3XW�����,�+ݳ���ʺJ)�'����e�{z����C����P���t/K���Q��������~�:��
U寪��^E��c��4�l�P�;Xgs�����ְ�\�&?/�t��I`�t;>f���s4�cz3Br%wЬ������QV2c�$T�$�����NםCKM��x��ȫ�Mޫn����Rm���n�<�:X�@���/�L���r���Dkd\�hT�FB�p����"s�6 Z����}3Y��R��j�<Qـ�������ρxڨy�W�C�>+�E(l�\-��"�D"��k�Ir/�+E��}�	"3��M_�7P�ݔ1�	��	&Cz�߾$P��^�62z���xȵ��/D ͧo�d}�d�4�uyV>z&v�%3��:!��t�l͔ä���Td�sR)G�l[W���bF]:��O���Ў�L� 0Q��2�6ti���D �q�ُ.�������(�����Ŷ�XZ�L��aX�z�|AV㩲�4w�q�@��ƭ�l��¥}'��~��i���D'���A֟�i>��l��<��U��[��cK� �,�1؉;O��r���+�����0!�lOƇ���F�R���d�k�T?���jIEK���OC�a8�H�
6S���]�b(x[-Hx���Zl9�������D��t����-����ZjQ5͏�U�zjuOUr\i��1�H����U��/	��	u��ʿ��݅#��f{�J��dY����J ~qËuFT�.f4#K����C<t|,�� ������7� �h|��7|�q5>��%~��IX��j��e3��6#��0��+�2�`)��i���l��i���GL�Z��cV7�~.�!k\�B�X�4�����S�4����
D]�"Zfm������zڲ�4s?��L��9R*��=\+�{o�͍��NԈp���Á����4�rk:@�/�m�1+�8@Z�J���%:]��m��u%ݹ:�f�J���P,�g��w�����?��/8��
$��/�ВC*s�vI}ޯr��m)���J��w�a�e}.��=�?���(ܗL�4�� VZ���y�+oLH �76� y�jqzv6�?�e�y���"��ӂ4��ܭ��uɛeR�����ʅ�c�}T#{پ���'� Ӟ���H�)�T�}��B8��)�e�B�5�v��/�U48ca�6�ue����l��_N����F�n9d�t�K \�-8�:��lܤ��!c�G���p#�Un9���&�A
����j=�������� ���9�F�$����g�б)�}�]���(��7�m�^�p3ت����:�Q����3��Ǭ�r	8̒�J��dpfSV�ҲJv����/f�3^Y�rq2� 9�)��εÁj��ͨF�X�D�xg�x�^Ѣ!*5P���&��f�8A��JSȟc���h��y�*v~E+y�o�Nz�����z����QVg*�7��]�Ku��
��	giii�k��iv��7_"d�9Kq�+��Q<Ԟ�}]
Y'm`�S�X�llLj?&��lq!�%ߡv�F�ū��7�6����66��p�z�Wd�⺸�_�c�2F�61���C�����\��ѯ1pCg���q��]Lx�b�׊��y�RDR/qa��NI��]H# PV^k�7���Bb��,���t�����2Q�|}��Q�����5&���$j��R��4�x�h���.�^�"ۙ����DJ�?K��&>������7�,ٓ�h\Q9��"��b�&�i���|���)��<*esL?b��t�����M��t7�س�D]R"%^$�����u$[泐1w9���YcJJJZ��X�.��n���C�S*
J���᫩��I�u�U�����Wڢ;�����DX/�Fk�rat��n�g�z/��{�~�t�*>��NFf�"�.�����B�\�jZ�1l�#냳oT�_t��ĥ��j?� �vM^_���`�u�	E�H��n���u�i�=���X�0��E��9k�}���i�h�*?�3�#������s�L��x�N��U�<�>C(��U�eV�e3X�[a��O�b�Ⱥ��l��}h�q���l�����D��W�S
T���GվsS��]��+Qn��/�<�p�5�Y=�g
E��sM� ���vm�h0�)Zs�t\N��5�@��K_���kV��_�w{����X�}ץc���7V��cV�b7��2?���,����Wc(��*6�j��^5���C���6`�[����=`� |�	��z�D�}c�6�����ٖTLt�����]��<��Cm�Ƚ��ݟ�,��RL��b�doTc�C�i� J����b�(G(_-�p)���͑t#A�ߓ�W���s�Ϲ5�6�޺�E�����dm|{��E�U�.+��&4�3�\ �f�	����Ⱥ"O�P�%�:D��,u_����E��e�|��2Y�
]G)�7#�H�+�>k�= B�-�����gU��շ�BFm��kױ!`af�wsy�����9�poL(��K2��lݪ�c��M� I���؛Sꥇ���$��
�}��q��움]�b5�,Vd��O��)||%###^$w��;*v��cT=�(�4>P��hP�P�m[��h��Jv�>g����[��tq�Zi&���c�W-�iR���
�$ҽÖ��]�b�
�
�,������5(>OMAD��-�ck��qt�Z<��f��������.��O��By��8�A"�6�:)�?��w�>���wz��z�O������~"�d�J�u.��������'թ�n��谏`�qJw3���_�A��I�>�~�mBCH�ɽYEP�,Tr���]ѐI��>��7�ma��%�����<�d�z�_!lT��Sseh��͒��,l�h66>q�$V�f[�� o�nGm/qQ������]�tw�����
?�V�<��� ɕ����@/c^�q������P��t���z�k6W��9�?�oovC�CGϐ�Y�7�(�z�hL�W�h��&qy���=����=����>�6�,��_?Md���#Z!�S!����5�Nf˟�G��q�Ad�x�
>|�>���@/��o��/v��6��I��^��m�-��ԈVm�	q;Sn�o�e���K���d���4�X�~��#���)���]��#� �ˎ�8�Rko�9�W	�b���i�\cΓ����KY��~�N�D���c3��H���41k��y��P��NZ�r���!��m&×N�2��J����Dm����B�m)1�o/����3�^[��Ϩ�?$��?w��m̕@j��΂s�f��{k�U��n�M��y٪��X^�F,��'̸�0E�AW�~[�˱�LdM}�����5b�O6z �AJ7�V<nVS��5���K���������n���w��M~�|�o�˳&u������ժFX�@v*� �|δ2��Pwl@��X��y}�j�(�_F����+�$�
)���P��E���� �)د	^f��(d�zp���a"sJZ�;H@������%q� ^��~T�̴k��)�t+�uI��5A����smΨx=�Rl�(D�� :�1jU䡴��0I�
ko���Zu�<"�L%?xV9�z���7��B;�܋�P'I��جZ�����UZC�uEͨr�����Χ6���mkc���^A���c���6�sRo�=��mE^�HT�4\���͠@�G�?�ޢ���oV3p�����L�&dKK��aI��P��R���Y\d�Y+�W��D��LF��hy�`� {W����wq��1�%@sp`��黛�2��[��UwSpu2�s��.��/�9�,)yy��S�m���W���/��.�SZ)%��~P,�[G����d�5���!�ߍ����?�V+�_^�i'��y��Y�6��?�ߥJ �+�� �3�Yorp�!Ⴢb`��4纾�e�*/%K�kҏվ���ZӽY���O"�"o�F�9��B
�;��_Wԛ-�)�?���$RZ�.�n�4򷌌�,'w��B�E�/���/�B8��bͨO��H����$���(#>oln��Xw7�2�A�{�){�����5�2���gCnN��K������ ��� �3��h�u�*�Bdy̟�1�&����8[2"���`�稦����|b�f�²�ⶤj��i��j�ÙN��_:<f)��|PPЁ��L?i�׻�w�Dg(��fި�Y�?xT&��*x����fi��2�^?�
u�����0�_A�F]�q8��#E(lg)�����v��Ry��M�g���Ǔ��c���H���UPQ�B�u��0��ݎ ������dV)��;eQ^�S)|�g���[&Fk��u��us�ß��8O��b��D�]޽sx���o�Ҙ���j���2��/�-�ٿ����s$<�H����i�!����Ki�\ 
��}i�Ł%�@���Ë$�ۯ�����O7��L��*zw�O����ס��'q4D���$1ā����S�uj��s9F���Q?�g����+��}=Z�[MA*��WN$��0�Bm8�ex��P���W��ۖ^.0����<���X��g�Մ{SƆ�n�Z)�=a�c���Y������R���lh۠�:���[�ڃ�C*�i�!a�Fłr]�A%���R��oVX��x��/�>Y#/��~0�4�H_C���7�:����ٝ�$d!��..ˑ؛䁥��=<{��]��׫a��-�����>�o6s�5ro㬟�G��T�R���*K��G
J�h�;1Đ������"l���9�V������F�B�� Z-vG^������yI���7�GZ�Mx�7;���q
��I�+�`�P,L��J�4f(�?���b&���;.3���Ѯ��W��@φ����pg'�!}��m��ߍf`ApЕR\[X���mӝ���̈́_�n��@*���j�T��DK�!wk[�3:`���Jʮe�N${�p{dmg�q!�q��m�șo�!0J(�vx)3���4������[��l
.顨6���.1!�7I�V��R��8�9�_��M_jjͷ��?��3����{oѓH-z���#A���E�DD���^G�ޢ������{}g�������>g���>{��hM}�nY�0酜�� ��Q��������eK����6��G���	���K
���Q��#���Ir�'�7��?+��`C��c*�}���ԟxz� v4g�KE�&���k��q���UW��q�{���_�ld���w�%2�p�S�>��{X�xA:Mڛ���2V\�]�ꖕ�{0	<1y��o�yz������	Q���6F��r}����u�8Ib���b��م�����9�Y��0_>�鿪��*h}��lh��
v՝���{�a�حƃ�J��8lsL� �A�W�H�8�LM(�F���$�����J�`MQhN*�����ɉkso��RS_/��9ѹ+w���5�����K񼽪�C���_��_��[�P�e'�e�餳�f�����LD{�\o������Ǉ����V3��Z�H�o�>��ײQ!ڶA)<` �ŏ��ɶ��e.�����ן���D���IvK֋��p�ɑ�x)A�/�Zin���m�'ci2����S<��ñ���z��MS>�#q���#ҝEz�p��[���y�r�`�"/dL�8�N���,����n/�t�ղc�/K��zP�����o%��:��x�j�%؍� �V�̠a"��;��K]T7�Aᦱ�;b������P������dY'-L�w�@[:&�����&%��+�V�fZ�'�?�J�z��ٳrM��[���){�Lju|/����K�3\���Nd����R��|�1
��a"�z׀�J ��Ճs"K`m�2���G}���_�䴡ɔX7�*����������������h\����qR �)�/�p�|;r�o��tص�e�ӱɃ����֛�}S���JFi����w�����<?M���-�X�H&]�b棉�.��͐�>���Z.�)�VU�z�N����$�MA��bykC�!���@xN!��E���f�9���4�҂z�rJK����1������;H�e|��&�/�E�ȏ��:��ೳO�<i��ߨ����ӣ<::z]C�C�TPP�<ۥ/.)Y�9;;yw{u�,�E�,���J���#x9R�UY�R�&A�����&<{Ϧ��~G�4�:��J(��ۡi]����0�_Z������|�_��;W�6-���x,�8�8�T����w١׫m915�o2��5o(��F!'%�˼4�A��9�h�q�3^��)횭pt�턲�ؘ�D�����ls��QNlu���!��$D ��k������ ���6ʒ...����[��=N--�Q*3y�� ^���Da!���(ZR�y~͉z�?\@(~���^�fg'��{/TBb�	+�B�*Vf�p?4�ef`�w� ����n�g�ms��g=J�sx|�GDJ����ʿ�ޚ��-���8���%3[�ɯ종�����{$%$F����y���x����y�I��B5�_y/�F����`pBb������~O��^�/t��+�u�10D��奲��i�����^	�9�3$����hu8XW��S��j��X_s6E󇗻w�F�G���kdX���"'N&7�(�׸�n#�$>s�� ,;���|;@c
'٢����`s8s-��gr�3���^N�Bܾ���~L����k�:Ȼ�k�:C�*�Tɩ�6M�}�<ݍ�	�9����11�h���6�|��SMъ3.RM,�$,8rd�F]��6:@`q�b�����n)�*�8�6<�+Y�7u�7u��я�U���g}䎈�.Dsd�O7e��/ ��3����4��mz�m����߸�^������{ ��Zh�|K�u(ޗ˔�J�� E�$)�(��ǵ�Pg���ǿ4�����n��NHBW�=,��k�����Q��T~g����r5Vr#uKR��3?"N�ʶ+j�氧ɨ1*!>���x*>U��jgdW�}�����J�r}�,ٚaV#"j�{Je>{~<;1�jA��H�b.�<Uf�Fn`b�(���\);��2���6��K^K+�y�De4ۏ;V�|���8���9F�4���ϣ�	ƧD�>�*}��S+]3����~mu���ĕP��\�����󾤤���­NmzBB*���F�b�݁�ZZZ��E�s���?�v�B�b����7����yF�B��T����D�M^�	t)
�t�E�.
˰��+"nϾb�2����`�7��K�;S�!X�}����0\���u�{aZg�{tɸi���]�x�}c�wXi�����@c��ø�'C��*󋺃/ͺ�����5x{�	`�H�<id���7�pm���KeTB6
�#֡�6��;l�b���[��H�Jy����&��.���š��''W���> ��k���#~�q.�=̬�U�Q���[m�9��=��'~Y���[��k��D��*�^д�qՊ����e��
Z�3xun�2]i��������S�X��|�w�_��o	��a\�DX�X�%$�n��M�*M��.�ɷ��V���ř�ô.L"�F�	i����x�Z�1���V�m��떇�~r�
O�-I��!&��w�^��={g��=�������#��f���QVW~iB[�;����V-�kg�:靿UL%���AV<�P�_����rs[�a��G)�~����V ��mp�Lq
��ފ��v����N�w��K�t����U.���u~�wH����dSq����,5[=W�hM	�[�������mO � �Q_R�_�@�gs�w]��ԃf#�sw����J������f/15<�?�.&�uc}y�.�� ��NqI~��0�P�c����ٞ��2�S�G� h�AD̊�N�;`������mvC�$������g�˔����|L���D8w������;��b�diGH�N����*�\��K,ܴo:H�ј�^;3���6h��K�g
�C?��u�֨`cUz�jH/��W�oV��+q�A��*�s�tp�TQL#j2�D���̺VfD�B��k�<������W
 ~W�����.1I�T|���F<z�yMb���	�y~ն�C'��뫊�����s/���S����IB�]0�;[8q<��q�FGE��-� �ڽ��
�HL3酩aS]�Y�WߟvA~�6[QZ0�-EO�ƍ��s�c�T�"����s�uT�����)<��'BXm��6����f83.�	�Em`�j�h6�3�c�˭�����_F��/�z���vgy#�	˳ù�_�{�B��/����Y.ꤟe=�	28�=��貓��`�T� ��~��&JT˨`3H�}u�;��η��Q�E��@�zv>�4

S�NK~��Ws`�b���1��ҹ;(���#г�8�$�|�e�0y����&�*�|�'��G4�q��:�Vi=����I.7���/�qŶ	ևZib&����OV<A<w��)t��Y��[_���FD���yH8x}�4BDR�S";P�"n��;���G��X�!��(�:�3͕�(��o���&O'4`O� �;�^s8����uv$l�:�Ď��D�gy�v�����"رԅ�Y�W�i�`���1�����B��|�͟��|��FU�kjz'�^c]T����w�\���?�:�||����k\e
��}�(����T��뇽c�7V�վxϣUU�m�L�x���`Lpv���U_q 7�6b��W�����_<��	)��[�u�����п�-�������{1O��A^�����O�Ž=u��#��?��Q�Q��R�x&ɄZ:��+�Lsh��L�\Z�'��7���Ik|�U���)ڣ�ذ���f��$�^��i21g��Z'�#��������׀���>W�s�7km�A��ѡ�8R�O�D�o7�bv>bk&=A�|I��"�<�m �u&0�랡�o��nu����:�f�KZ��xEX���{��
Q��a�m����C�-�t;�e=EV��B��/Q�ᔐ��8^��g��Sşp^�މ��t�����R�bO�t�ssv��!	{�Z'Y����06jc�q;��.��Aeo����w�d��k���.�:�[�Cm�3�Q	}����-m2ch�n��߶��%�\��?F&~��L>|\�����f��[����3�+"�����(Z��_��Ŏ�	�=M1b�\�/^�(�u����R�2�YvnK�|+�g�T��n�B$��x��H&g����h% h`��D��ﶷNN,�"���`?-��N�b���y-�t�.,��s��}��H`�%����&��ٮ�3��?e�_��͒B< �}7�����; �g&qN	�b�G0��=m	��Y�������q֨�~ei�7bIE9k���'k�F�������P➳���Ew��HD��j&Kxx� ��2ݚ�8�/{��5#A�߰�y+]���y���I��3�}��/�l��F�� �$D�O~���W���J��%�&�?H��Ox���I7��,��+NɿJ� �#Kd�����D�����*j����d��rE��A��	�Z/�}��H0Z#P��3,>��7��DK����_r��,���9�d�L�p��X]_�J�i�ãP<�q\��s�~��S�m)\��Yij:�}rIPyDр�f�����S����{�2�S�$�NZ�Qڡg@@�"/�Ct]�d��t�V5�Gڜ)�i��Հ� Zw��n�z�����q*=3.P-��\���`��W=���,o}�`�6���������"*�_s'�t�2"�y:4�b6r�ik��Ͱ��S!�Ѐ��	�ah屵���Q�cQ���4���]G���!��	�\�%�Q���p�O�J��?/�'�-S�vuay9�*��6<҇�n���!	�d�������9w�&�wJO|Y�$�bw�a�(�y��H-�����|bp7s����@����*X���R{������Y~y6>zĚ Vǳ����F������Y�ɿ� =�(���Qg\�m��Q!+�xDb5v���x��^ ��J��&���j �jqK�fSƿ��yC3(�؁8�Jz6�̕et�_s;���"�7!�uT��C�!6�~�{1��j�H1�����[��;`탬7t?~�>�z8�aq�{u�7� �o�����Õ�f!T�Q��_�R$�<�*�u�z�W����/�N���)��z������Y��&���M��X��3�P�">��0e]�+���00�����M������6/ND�����B%��h��I�d��`��µw�C����s9��X5�B�Z����~7���?����6.`����_��"�1���n�6~�����\�Ĩ�&$�?�U�M����Nj��CAf)�%��r�z{��0��%��ׄt�2���I3.,,EJe56�P��At-��F��4�&gg<����Ʒ���²�EΧ�I��<� �(h�	��$k�sB�)�=$~#���0���7�9�/�q,+�c9��ʹ�U�.��/��E�S��0�P4wa���n��mFU�m�b�>9n�ց���ި�@a�����(�P�X�l9��JQ�B�2WJ&�������L�H�>�ϐ��]F-�9�{�ɾVR�?:>�w���s� ���r!�|:�aS����d��s�rR���S��I�Q_�L�yc�)M��i��n�6f#iqȘ��ܙ�bO_���2�����ȟy�8��V������s��fۤ^�|��Q_����*3�
۳��8���6#�Gl�Q��t�����ŧʋ�:�:�@\(��RS_�s�%+S0�+Z�B-�Z-�d�b���\#eggg%�o�[O�ߖ��&�LG��$A�G����P䯞mb���23GJ�*K�ﶟ2�l7���	qq7r�Q�[��mMz�~ �?�J���W[�"�X1rL��6%㰔V�n�����c3�=!V�����t�(��.�T�P����uض,�D��6�a,H2� �������vG7t�ƒ�M���ݙ���ȨH�5�v	ʝ0���zT7D�a�K��L�SpGQ>�D�eJ������ ��(�p��1e�9�>��b�N�N�z�N������I!�3c�/zb�<������V��VPٞ2�������b�����5�k����@d_<���N��^GlƿvHRB���#E�Nr��:E	�$�ϟsw�iDO�kp�A�L��±�'W敮����֘�=��;���jHNN-�d���D.�j<e`B�8��ۡ<g����>�/���V�a�q�
��}����FF��O���A�^T��{��Xg�'��#Z�}+��|E�m7�ݧVkE(�YG�2S���'7�SC�.S��j%��^�u�[��<��;MJ��A��rr["�Q�u&	 ��G�;��|�;'���s��Ѥ�E��D�����Y��؏�w��O��o����g�G�֢m�D����W(x=���o�e�JӊǙ�������A+}_s�4G�ʁ��D��OH�JɋBŐ����M�x3{��*��}ʇ�b]36�Y�D�C稼OTm�-\]u�
9J1ҞK�����=��l�����ޟk��O��G�}b21�#d��Ɵ�R����KO�o
������Q�m-�����M9/��l�|:P��ނ��݃?<��q�VB�RPT|��>���~۟u <�"����ayE�n��2�G�~�7U�^b��p�s����xr�E�sw8	�����?��ԉ���_F1�����T^ؙNT����^���:�j�p�l*A��o���;pK��("�ݍ�w��i?x3��F4brfU���0�1�ƈ�o�ؒ�� �*Ҭ�b*��Rp�03{�k0={z���%WA󆳺��톂��L�����Ǭ�h�i�Cj�H�M�fǩ��$�t�l�lϐ��ypu�=��d$�ӱ������5�x��Z�4���8���4���AZ��dlޯ�%���Վ%{��&R?��U��o���x�B�)�@(8~T��
����'+}�P��� �AVzZ(�,���_�A!Yx*A��]��d%̹SvOP�[��A�x��k�O�)���@�pLL���LS�u���W�6��im���������G��C &��9���YE}/]�o.$BAj4E�y�Q	�6�2U7-�a�sk�2R��P��fIYV���EW ����wzQЛ�����6����i�䯏��&�D��֩'d��
ˣ�F�P�#W�Zɦ���'Ϗ��y��rG�@0^"RR�XN]ug;����-�.:E��'x6��Bg���{P	����V�y���=���]�k�~�i���Aibrk'��1:n&ߧ��YS�):ByYg�҇�?[=l�A��"�5���!0k
�{�����o��H�[qiq������ɷɩBڃ!������.�.���R�u�X���
�:�f�ĢQl
�� ��Q:��\��[	H�Z�����}	��趤|�P<!�/R+$G�czT�j�>JIύ�B����@�dI�.�ܦ�&���xkC1rw߽]-���]�4Aġ܊��|Yv�0����y֩NX��b*�`��<�x��	��>~�ɧB����$,*�r�܉����ú��ۗ8��O�ASL��s����Z}1k�F���t�ǿw�~KD��t���,nU�[-�c�Iԕ���G�|w7��I�+J���i#�&��5JH�5s��?4���nJQt��uqq����9�T��Nf��C��Ӳ?r/D>�V-�E�Ț%��d�N�3�C�� A��~��yFp�A��9��>f�,kEC.^xA����S�ݩ�&�0�i{�r\�x���ZX���) ��Y�!<�1=	A�s������^)f��u�Y2�K�p��Z�bl�������gB-�sr����!Q{Я^��ޫ?�P�L�'�[;�v��1>P�ѣl��л��Q�αv`���&���7؉���˱�{¶L=�r���zG�ϟ??�?W78��7�<�$����	�gY�\�qss�]ិW�Z��C�E앒��������F�ɣ/����,أ�G��t�Q� ��9i
V���\����C1��A^�k�$s�	QN���,n�Aq"ߖOEc� �k�1w'�@�
ӓ��d� �x�A<��mu=Z��ˈ�A�����:uvO��B��hZ?�:ԝ����m�Bg��;�}̄ǒ�Y{p�S�W6��:���N����4�ߢ>[���QbX�45�KXOZr;M���.U(.VT��K.�z�/t�0�`�@mO$����i�P]Z%��YM����6vQ�te�[e��)!�j+��O��gE��uII��]�/f�=]���9%!&�@9�Z�\͉>��*J!J�za����m(]�r���2B(yG?��c���6V^H��GBˤ(��yp����J���h�/��K�
Ry�!�5�Pv�tb>�R�O�YP��+�qm�,�!��Q�ns��/��I�:��K�n����;�O��~��7�̞m�B,A��"�}GPIU����8�@x^�o!�M�2���2r&&���('���Ŷ��R��'$t2��n����Q�8�i5��B9�)�i��@��(���+7���h�y\JHNOO�@�iT���9�`�\�\�/jӡo("��~�����k��2�����;�o��^?��8�A1�� �hv���w�vr��L��أr��_Rf)Tfv��"����]aP|������@ ��>���y�6��q�5E����[J��z0����o�z��H�/k�cG�P*�cN�p���ÏF�2{�0���5*����z���x��8!�O����xpᅻ&���3...J ϲ���>O�16xB8F�lO{��;$���o�#f�����ΨSk���.��Oz,R����������n�u�;�y����(3�-,@�bY�؏陙{ �:iF_�
��kQ&�E �X�ޛ�n�3�<�IR��"f�i�^���}�V��_��e�(�ZJ�	}Fʕ(�ѥ]�q���A�Z
���˸��QZ'Պ����7*�����l
. #�CAx���H���}�`W]�G�����O�
���ԝK����ҹ&��� �NO�'^�}��x4Y�n�B�syP����ҌVηF�=�q��ۛ�ڦ8�ߛ����l��_tL�F�L2��_n�����5?��`������4C��E-��y���l�껐u@�zt�r�O�b��F�i���Y� �����F�3-7{Z�����\	f���U��pv�_|,
�y�g�<�B~O���q����uH%x���\�Ȧ���*�ל�ڐ��Lby��U������k >%'o4"onz`�n5[;_�n^�0�L�uyyt�8���ߛ�����=IpR�j�K�(�ʮ������!25��R򍅩���h�>d����1i5R&�ht����7��7l�ZG�'�S���pjg,%h�8ǰ��6+	������ag����V�9;p�Y��Ly��,�����ݓ����,�Y�#�a`d<<ZS��	��P6�nL�e�e}L�>#�Û���p3G~G���Q�*6��+0�2(�D3�i����F�0�<k��<y�,�$� �X�呣�j�#�"���ޫ_j�T���K_�#p/6�ŻM �{n�݁{X#$����?�ﱏ^9:�Ⱥ+��r?��OD�ٟ������=��I��8dؖ�ާ?<7���>K]
�۝���z��7Ω�f�2�\{]��YK�c�� ��i���A¶y>L�ub�%�M�1VQnh��.Щ�DW������R��g&��-���>�z��5K$����qa���FIF�����j�_�<Jc��,�aN/���p���1��E��~O�a\3hO��D*��J�[��t6���>��L��V���p֚��Q���g��lR������X���]�m-����c�j�3���lw&x��nP����I���Ѫ�?�����_�u���k;�(%Y�����sbs�7r8Q���t ��P��B�զ���c<t���PҪ�ož�*,N����)����n��`�A�*���%)���3�)*KVr�E�h��W�\�=bz�h㽥��!HK��3���%��@)
1�u�wWz[E
X�L���8�&Ys#�1%uT���Z�˞��-G�5��|�5+�k�7�=#O�V�5«+_+�Szn����t�$WnG�<��Ep��V��D�;�T������7�3��U��J�C;ִ�/B��{@�����ܢ�vL���0�S���u�^�%}h@i�Tpy�S(
���$������
E�Ũ/��<- SR����f�qK)j/����/�T��Y���+*#�0��C��0e}ߴWs4u�(�s�&��B���Ɗ�єV;s��ot]l��(f�����z_m�-T�3]e���B�B�,�	7j�@��̀3**.����@��`d����� ����2.�Mǰ���>��6(�=�1Y�5!y:;�O>8�P~K������k��Q��@v����T��9���^%�z�-��4xY%��:� ��c<��ᑛ46��!c�;*�V���[��J���7>��ދ�ܿ��2w���h���u��7EGfS�IU�,���	u�t��?[8��<�b�zs���Z��p?~Y�jc#37/s�&ݘK�����ڴ"OZ<���C��q%�6x§s���5���{�
+��qI'�凞TVLD�'"b�nGF���g���\(�1X�Q�p�����,hS(���u�Л�P�*���[Z�hm}�CU@��-�^�Dڮ��ݓȋl��ǘreؤ"@���Y�r�������gi����.�(����}�G03����S��A���)t}�#��\��N}$����qd��5sz\[�����K	���Y�~�dU3b^G�� ���{?^]W�X�3���x����b@�;�k��J��&d@+F��$�#���&�C���� _�@�0u��8"P��ٷ�?���'�*�#`#��L&��	�ΪA6J�9� H�ğX��2���MYږvO$B�Y�'2�.C�;��Q:Uܣ���?pFm�d�h��ɗ��\���X�o�����p�!"��&Xwn�����&˹�Y%�0�`��)G9!X�h��C�[���_L�R�,�Гף��n}S'I��(�D�P�e�M[��]�e��:�5�����`R%D�cgVN�������Y{-pr��<�WC��sd?2�E���H�l�'���w�����c��:��^��fӺ1����y���p-9ߔd���D�z5�7�jQ&//V▩Ǧf��|U��9��Ƚ4`�ӗ�b����[o�S�������M����-s�[,WX����$��1\�!sz?��\�؅�Q�ϟw��"S���[
��u�9f��<g�8	��8r��r�ݖm�D����J�,b��%�+�v�8_Ё�}ű�ߓ���Н��Z�N��h�"*0:���ھ@�!�7�$;�:ǅ�H|c$�����r\����?��A���4N�E�&}nh�V7�>f���Z�̗L��� �C� 
�芧�FȪ�X�����c���'>���~��4~����M�X����#	p�c3õ���w���p%#Ƕ"7M�ьR������͐��x��j�]h}*��a4����l��P�}	�U/[����xS���12}��_�=��d��˧����1[�l.�5^+}�2�Q;�Ȅ��vl����:��׿�w�qϨ�z����ͪ�,�������;���X~K���T�R"l�_�OÓ�o�L���m_��9��b�v\�L�5�ҩ(� A�a���FU�{����\��O�N�=��p4&t�kK��N�%��Z!B��&VP�����tx��"�,��|���ʼ�m]�+��7�:�@�����C���u�oR��PvOZ����+� ��(��F���"U
� 8�)8/w� n��:lZ��	��VwJ�Mu��tY�mf�o���"�:I5]?�p-���H�E��g���eyK;S�w�x�SN�����^9���~���Go��A���b�����>zm����I0Y ���冿�H2%���M*�Ŏ���G����(�lOk���?`��"fu�8\�E��w?��t��c,�}w��A`�&1�&���\�~�G�r/����H�4!f t�4�H˒R��}@&q����ݎ�.�C�<f�ߕ])���(|1�	�1�$���8��2mq�s�}S��5F�J����V �U��m�����?��~oetmm������� �60��I�9'Z`\`����{κ"��{~���[��N�S��[ y����yI��U��!stK�����#)���Y�$��)�(.� ���%��*dF�\���2��'Ŧ��o�޿�0���!H-&��dڋ��Z]���`$J��_8��22�tiL�T|��_�_������ݥ��7�,n�o�Ϣ�� c�� ���ȸ�����'䖎�+Wq�A��}씰��?T�%^V�E���Vi8�w���ʠ${����]� �Tq-k��6{��1Kf(o���jOk�aaM��Hy͛m%���T�7�Ӻ�[pGa�����b�8G���}�o��XX�|�ú�+c�+�Bfy�>��N1��5O�,e<�%��hn��^7]�8z��x�2� [���x���T���oy.�K�|y4������Ϙ�.��]b-W�S� %]�do�g9V�{����N1�����Q2|e��3o������%� �7BXs	s~D�vy`��^���إ�Ҳ�e��ܘ3�{F�>���/��>=Yߜ%y����%=��Z �ƌ�=&����I�ܽ4����[����(��#'N3ÖK��ѣ���r��?�!���O��3�6̘2"�Cep��/�I	x�qvGv&�����K�犜��Z�� A�����^R析��t2�l��]�f�݇W���Y�{z���*�>YA�jΏ�~�V�o�lk5ӸO@�m�&���~k��g��/��f�SU�[aC=�~�o�'����k_��,�0UiҞv�o
�%e{�-b���W�k9E0��l7�9H���E�o��dR7�Z�@��9����w���(�&)�ft��P�����'���Fe�N�<i������1l��*D��MM��W�,�Nx33^d�4 ��[�6l[�l���ħdsqL��w~���f����'Wo��苆Z�N�&��,���$PH��^��ͻ�<���Ր���/#�R�0#����X�G9�ԫW�m�ug�4r0C�y[O��F4����4�9s�%�,����2Vh��I�t�����:�A���[_q�y����Gd:w?yG� >gA�d��v�Cw��! G�	<'U��:J�/Ѓ&)q�Ò�l|Y��mV6��T���~���yt��y������
	E�`└��Sb�FS-��T0g�M`���c�c��&���v�w.��,����b���̴�.�Ż<�_��S�`�?�C��k.A��Ϟ��
��B	��cIᘙ-��.��Zy	¹�f$����}�=��e��[����Ãe��÷UUU�����7���!242J��lq�hn�Ӻ���ly�`�9�?�a����y��筨�����"��b�����90�����J��[�7��������[1������y��@Rn�*��0�(|�z�/�i��LE�&�h_m�O�>:j�h6W�3=3}{Gǃ��Tn\�Sޤ����u����9����u�9|�|qd�|4�Z�!��z�[�=�y�kr�[���]ћT�?ۆ�����;��B���5��JI �d�
�=�7m�C&�!����＼�g>�揿�I$5Rb�/�y�����u���'o�!�n��q�|A�r��	o_�☲`n�880{[�'�o)+#��<��o�_�Ei	G;���n��}_i��q%x������ԃ��_v�x|y���G��K��Y�V$�f|�[��Q�u����v��ʔ�Ge����_�DCK���c��ż$���jlj�éc��H}���Я�׫����{����o=��yX��X(��{]\[]<F�w������SG����F*6�܋��[�~8CC/*QLW��m_aʥx�o�Bg!x����"?�����SR�H�oRgG������K����,�e��/*���;L����F����ˑ%���)K�<*���R�o�>��j��lo�V���Io��IYt�xp%f�ڴ '{#�%�"d��#JE-�5Jv܇\C�8y� ������D$�9y-��|J�����D�OG$E��n.�J���VzY��67mm5��6��SS;GG�&���]��.���1P� ����K%5�P�g���yg��QW'RS_o����R^Z�ty�1��Z�x�)�@��P������.��8A9 ����wB3�xg���A�|ځ �p��W���Ʊr��֮�Q�瞔�5�ߚ&�h9�!�E=P���vg�~_8]~�3�Ǽ23Q�y���n�!�ڧ1���y����$:&&�=C#�{���
�&�6�_G��>&l�M����{�p5=����v�j��z�[�g�&��Q�wr�(���aPe�����b�%܋!�T�KQO�0G�Ƥ�`���^v�Q��;G.C�c�y_��na��3<=g{�������TS=�444j�k"��PY�B�¬�p�����:��{�T9���p�o&-_?
�O��֖�I��k����o��˟��1?-H��1�ܷ�ߍ�2N����l��^��������%$V[DSK�d����|���"έI�9�?��Ӣ�iZ��W�E4�?+��'p3�y�[4�N�����»0J�j*����ɔ�O��{�z�I.T_Gcch�e�Z:7�v 5q�MGs#Ύ��DWـ�_eA5�z�7�f����Wv�%�8�(
�ׂ���t#�v4|}��(?(p���XA�-���>8]��ޜ�����>kY|M��m�<m��#m$���4�{�,^Y�̔��eE�sg��p�ͯ���{�����V#�sI7��7,�S'���Lہ΋��4��_e+/���H��_]�t�9�K�<g?+%|��\����Ua`1<ʯ
p0��9ğ�y�;��ʩO�*tǛ<88辣�8��;X�L4v��z��n��q�~v�K»i�C���$Zv�RS��P{rޏ]Yڿ[_D������'���[H�D��Q���G}���es����=z����676��2�fAߞ~�;�����!11ۼ��{�G������ȑ������:G�h㤠�!C�N6��W�^d|��֎���r{�//�܁555��ՁD��0�
���P��H
G��pi�pm��m�Rs�-��#QQ�bi��0�g������v���}�⠼�L��Y�-)�́��X�:N��ꣾe���*@�Q�'	�t)y:m�Zdü	m;�J)�b��U��g�jȪ��*��)W���-���?ƅ�� #Ejs�gz��j�����6�2��.���|�����G�B�p3�˭7�|��������//-$��`�"�u��|�)�n�,�]ˍ���G�PG�9�,��X;&���|݌�<ވ���2����ν��0L�R�2OW#& �ss���j`oَ��/��e��_:[��.��i%�z����������-��n����{\�ܭx��˸�G�ߪ�5�T���gf�����#c�Zh��z��S��keg׏v�U���]1%����>0W�ӗ�s���`5�j�*9�Ih)��^�[��|RdZG@���	��j��ׇ`���5&g~��^��[��u��X+��6�.D`�j�NlM4��6����H�O��P4�I0�+�a�.)TX�{22E���ھ�8��,sNJoI�,�W�|�w>� o}�X��i�Wo�+|i��H��k��5����!�<?�0��ͧr0 �d�e�06��	w:0@EM5�������|:p<��〮2�09������4 �[��B��P��V�ǝ���@��]�紿��|fKۓ%E���J�|oFH^35P ��=�iqC�H�G����ސ�VJ�;�l
v�8?(	��k^��<���s�,U;���8����S����HZ�?k'I<��檅��~OzoN���
��%I��3h�qO]:|ll�B2��H�����fpa#��w�y���"9)��&�4%+,��x�t�lxU�ҹi�8���	җ#��C��Ȣ���]n`z(��?�mo�	ò�£*�	�P�+!DVU̓�����'a�$�±����"�bn�L���y����_�.�u�e��ޓyΆԅC�_��M)$��h���u^�!.��!0qM���LF�0�� �TS�)�z�sű5�Y�D�{�����F�k'�i�X���_��xć 6��rź/2�#m��쮞�a�!!}ǡ��M��ݪ�-��TH��Z��;�P+؈_���䶋�8Q��#�8QQ��ُ΁?a	b5�_��e	H6.��?u�ם#�Sp:n��u
�yo�ݻ����*8��E)HP������)�-����+�q��"��ri�����M&�ZC}vQһ��e�?�����S�Y�w�O|������?BN�O�Q��¹�$]Jٵ�f�/˥�����9��+s֕g���G�u�C���J([ȦP���EHFF8;��l���PvI%�y�93�Ȏㆽ��-�������p���y������~�^�.0�7��N7�t�TE����8��?�Yp��ޝ����~�IL��'���wg�ݛ/�Th܃邟�"}<��N��Ê_�M�b�H��\��m$Dw&N�>���t!�7Bk��G�]s�zo����DQw��D;tO�+�5$T�A��/�ۏw;���
�{n�k�.���!<b�m�584� �c9�) '�l���
K�����<*�k{<㩙c&X7@[N�8%w�5n���vi0���:�����C���oF��I�S�3=��{�+j�=��OD����t90���qp+m�X~��lA"���:�y��ݙ�!�sF��_*u{8��gu�*]W� aY�7|V�u�"�S7��CL���^�Q�O�>���,�~�'ާ��dgm�3�+�fVV�}.���O�);YӉ'ȿɀ3�;�wr�md	�̷cy$6���(��~oj�&���Ϙ8���|��.)kOK�m]�$KH2�Һ�nv.���i#���%��fb����srU$�i�R3o��~!��7���P�K�y�d��U�:zs���~���/R��v���:�X�A2�B�ٹ 2]">6��ٌ&bd|+W%�Jbbbq�˳ Kl@�T�{
�%ꅆ�Ʒ�P���_��`�*b�[?���(EQ1qm��[���R*�a-�~���<[&3qa�q�9H��m������s���;V �N��fu=��=o��3��%����1�ئh��LȊ�VB�b��I5�:�${(�*�{�ݫ��N$θ�q��+S�@���n�㌑Q�������j�/Z@��|.1,���.����-�y�F�3�H�����������mCE����dM�yܴ��7���Z�]�D<?��M��Z����e�JN�u��>6��(�ǻ��6ҊJ���Uq�g��oS���bb$��Q�]Vv��^OZJ*�7KB^bb8��}�e�3����ܣˑg^���SԤ39{��ki�o�_9B�B��8^>�j3淍2n�{����N��������m�Ý��t ���>�QB����_׆���SWpo^x�d�5fl� �"����#�̞_zd���&�;�Ւ�j@^ �9���ύ׀Y���"����򮠠�$������YV���W+�R����_��TUk>{�K�3z�U0�`�ڧ��6�f~�a�˾A$�W)��\T=������U���'�jc'L���]7V�A���}� ��%ր����`!V�h[���_�dq���Fɜ���z�r'��B�R�4�>�
��W3�1p#?�\W���rX��8h���P&�?��^K�����~�K?�7h|����D�nd�8��?e�cOR0#��2�����k�B�+�G{�uc���CJJI��	������������Z��>x�e�Qڕ��g�SOa��X6J���;����K,�9<���ҍ�߈b�x�������'(��ƷŁD���������T�mD��>){[�L����������w��{��&�F�/��R�;ż�iu�k�&����߉%;�w�siǮ�^�}Y��޹�}K+\��T2J ��IsU0ݴ9}v���e�fO����T��3+��Q=��X�0�2��5.� 6��Y�ҸM��q+� 7�*o�T���<Q�+�;e����`��?u��?L0�v�ػI��b�zy�dqu��C�%�.��>�/	=~'�T�6x[ǐKB�KU��Sv����[�q)�nzo����K|��m�8����R�`�̔��:` 1��I� V>�P�ȥ���:�| �d���Q1Z�2�u�2T�,99�,�-��l`��t*�"���t��~r���V��D���?Y2�:�^3��q��aQ]�I�Uy�?�F�{q���wl-�_s>:��V�_u����ڗ�0-�gϤ�u\&�(q87���R�H�rv~dd�?D�WJ�D�I~��΂�O� h�>�T�$uU�6�x�	/���� G-U��$�R~��z����<e����򹌆�
Z�'�n7�b5޿x�ٰS�@@��&m(AH�r [�{�� �3�9E!����B�E�_�1�wޑ���Β+r�8��`}tR7��͐v���`�o��Ԁ��t���G����tRi�8�#�(����t��ژ�J��')��.���:�
qzwy!q9z?o��C���O��'������D9�������>�����r�����T��Df�G:���s鹒ᱺ̱�Ci.���=H����xT^4�����,s..���-�k[%7�Vs��џ��L��ߕ�� �������t����6��HN��T��$�V�v�]o�ǡEX�#�R�]/0��GKMET�CV8�^�)|���|X��^�����xA��~G֣D�&� �.p��t	_�f؂��WVA�^���Є+�K�ܖU�i;^ի�1QSS_��P���#^��
e�_�jh�W0������l�z�`�h,+N'QV���V���';�n0����l
��~�f��V�#+r��3i�g��m�_�?L(��T�`�]t�j|/K�����z����r�Y���eF��f�l�gJ(����6�;;'gs��[�W;	4.�[7D�6�|���X����8zI�AȐ^���qo�N#���ys�ٞ�MT�퓿�x�C�xi@��ôz޽����ф��Q�X�Yէ�<J����F�?�����*�����j��W����Qɏj@O�p�
�	�\}1f��Q8�Q�r��ǩ���דy�)o�C�-�3�u��A�U��ؑRWO�e����č_�>��M�Pz�-w���ޕR��N�Z����Q�^�x�Xkֵ�|�]ҭ���,;/(y�+��������,������(�N��6�6�_��ɏY�eNI{���ֹ�+�(��y"l*l�"W5���$�fy�s��[��m�}��xA�����x¼��唶l��k�׹?;���+T����N>5��%���)O�l��g;F��5�x�u����[݋F�ͺ�	�T
�D˲m��uu_�wn&�QG�˅Gu�\�q���b���M���j'1��܁�YK��ҩ��'a�^��^G3.����������r��������A���2���eWq3F�/j@�V�����!�Q�^�����9	XA���QO?�-����X��bZ���U-��r�?.��{�=]f�)���sn^��k۫EGr&���M��<6l�4��kW)3+���ڇ��4�r�6��b��}� �;lY�yݻ���<�^T��^TkVҝG9:!bVL�?��V�-��K��v�`�ԍ��ŉ7)��}6i�J�@>�]5��c4�ː5���tw%fx�JD ��0BXb�N����V�I5tka���'ğ��\C�RG��ϡ�G��0�����/�[b��K����	'��\�R�����������D�,q��l�7o<C�3:+�X����2=�`�-��Gu��|��Pvx��t��(���x�]������⧟¾�4�J��|2��Y�o���T�#��/cK�?qy�s{�mA~�i���q�i{�;I�t�ƀGAn���>nE�����仩�o?��xM14�R�*ȽI�K��|V?U:.��O��8��3?k�}9�X�r�ܡ��K�t�?[�h�U>�~�bp�i�Q܇z�rq���n_��:B�G�M� ��=�B�&�b��f��.����QCp�G�Rr����@UC`�䶖�k)�KwJ3&sa�X3�]_z�y/$��7m�R��2�jd�)h���Ae��(~q̐=�w���|����پ� 0���a!��I���O�,t�j��SQsHTO�����E����|#g��1|=��������?UԱF�6,�x��|V��5�oWď�+�N{C�O ��"""��3��G�vI,\zO<�\��~N����+6����_����N�R*Gm&ښTJxtp�0�����������ALej��4��\��N�Vo���鄚�r\��fC�--�~�ao!m�u�m���JK[��� ���q���iJ�,���?�3<`rtr@⣗�C~[ZZJ ��W�V����&�u卦8���!���Z��@~L�[�]�;b�s4���n��ė0b��������NU�_r�8�+1����Q��\�5��X�kUp2���"�m�{b>�V"������p4k�?t��B�P��+դ�Dt�4n��`���(�Л��Q*Ȧ��ײ�A	\��p�@�������W�<���w�4���ͽ֌Pb�G��������S@$����k�垺K�u��[}Ɲ�i�&�u�3?������'����(��
�z~BOAZK�[)�"J��[xL��I���s�,i ������������T�����<U�ҋ��Ї��V����dϐ*r��&4;;�junD����Ld8\�jPB���v�A�+���u"|hA��gE������7Aao1�>Z��!�+>����L�f/)K�=v�!�AJ��O���,�W�p�T����`SV�b�R
�_>l�f�{��'?5M� i�����_�Ik��+�B9:����3�1���<�$8\�������=X�ͯ�����P�-�m�W-�D�6��@�g�<���𖯺c����?G�,��?%���V�"{Ž6̺#rQ��yq����(S�Χpé_bO4g����*OlC"8c��Q���!�j��;��1E��*��\h���[5B����L
�{���e��а�I���˾�*j���(:O�7�,��I*�{*�R �d����͏r��R�nk�e����4����	��QX�=�E{U��7��j��.��'����@/ؙ�K�Լk�"E��Z��
�;�G"w0�}1�0h�:V:!�a���c�_�&����cep�8��՛���2kh�[]___�T�a�Q�N��bl� ���h���i�q�о�m�:1��d��k�����[/2ֿ�`\���+�A��A(�M~�
D��j������
.��O��e�����Ԋ.8w��睇�!Q`�g/���ppe�G6����F[��6������m�6�Q��Pg�:��o==T$s��ML��.g�½!�7�:�	�M+x訾'oUxk�N���I�".�/O'm	ǣ��m��=�
_�]Ѫ�{o1�+H�~�V�Yո�[��z�:8��
���:�-�}[���+M�s�ᣛ��i*G�˓�;��Z�%w�����Y�-3'��~8 ���J��0\��ڞ�E�&� �KNu�8b"�����ٻj����eK�"��yߑ��;4�{�w�?�v�����684�F�q�9�e_v(<&��>�B����IY̛!p5<,��,˳i�=�#��o|{4 ��ZAu�jbw��N��$�����^�����G�T��h{�1	���I�UXt���G3:�Zj�[[���ђQ�cM^_�QTZ���TT�����j룇&-ˎ����{��U�ؕ-;����m�d�7��W��F�.��UA��.��͑�� ��D\ϾƠ�[:5=���  �Α��`e��w� ��C�o?zI�P��M�r�[��D��˦�۳�$��8w���Y���n@_h�rXIԓ�έ;ƃ��w26c�Ėdܤ������Q�+��Ӫ���_�D���-o��>� ���t������&.��``?��-�h�Zb��s-CԀ$�X:\��P'�\����#�|����D��)��zz�SU���j� ��`��t��i_���LF����8�G����߯q�s�;r�^yNP�ӸR� ���q��z�����mm<c��,_�Q����c�F{����y_>(�s�<����l̎'j����TҸ���&#>�a�I���C��^��~����r:S����[ uL��~A`F��		�z��7���U�Ŧg��7K��PP�����f��H�q�j��I@m
{�1���ۍ1���X���&�q�϶�$1��j���L�
������J���Ι��by0B[n��&��>�,�E"�>�4ݙ�6GCwg�tXϲ
�)=xÙ �X�e�Vt�����1�Kךm@��:�xVv.ޛ�#����������D�v�W[6� ?pj�%�v6.��žVdzS^s{�8�𫨷)�ŀ��);����Vt{ښe��e�W��T_1�,�D�Iɳ]ץ<�}�z�����1;��¦�T^u�C���w����J(|_n;���B����F�n�j����đC<�>)���G�u�W&#�2qlT��:
�ꁷ��\ݦu �kB��ҋ���q���mQf'��ٔ�'�5`�/�3��Հ�1����kx>'�����5���;0v¹]|��<�/&U��}�۶��:���]�������0�A�������y]�_���,G�=����D���6�����d�A�55u��B���Ə�+����m>|�pitq��cؚ]���1���GH�y���ε5���<�=E-�;�|���\��yb&��N�����tS��:�ӡa^\ǫy���[�9@�#}7�¶')��:���1��&�\�}z(*&����Q��\ɾ���cd�s&I���\ӯ� ��w�����&1��^y��;Ys��v=ֈ�ҹJH���?������F}��]Ϟ=�c�%a�I��FvvN%x`����ҭ��1p>wSVO��{Uu=�u!�Սj���%������iP���_��bjZls�B��(.G0�.�zU-Yx����{"r����]�Vlv0VN��y4����d^D5V�8�&���hz��tѵ"�c�_��c��
<���\8�4�>��3b������%OU���kmi����.�?�r�d�&���@6V]gy���v��g��F�~��@����l���V"�)4��gt�qoHws�D�i�L{�TM���#:�ڼo�ρ��z	lJ�[_熽h��7SݩҗSE�Ӥ�wf����[��x~���v��9�P^�`}S�jZ�hD�i���JF�E�C^����٤�����h^����*K�q[e^+v��߷E�!V֋���߸?NW��f�G�W�7q��gg\�dK���9��W���v�u�^׆�~�2�^c���OW�M3�lM�m�(�
�P�V64��E|r8􊮘��!��E�΍_K)L���b	�Xn���f����?#U5�Q11�"iR&%r%��>�,�m�nF�ش=sI��y{P�������CR���{ͨߒ�1/���P������8�j�G�k.�� �2;�U8���;nw��z������'��1�aP�P���#����)�kn���$>��(�rk%�r�鋆(�>}��5וL�3wV���;{�/c`�֥����� A-�{�ޛ~���ٕ��	��8���������ɔ� �[�qq�������^�;�m@�K⧭xK	j7`��q�\w�r�q��)Ks�-�Z���a1ٝӜޤf;7i������\�M��ĩ̴�L����q9o���6�m�<i}��_pSS���b���Y��~�'e7=w���^)y�ߜT;��h���
R&�=�/�d���D���߁�%�g#����F�T�������V��k�m2D�%�fQ�_%���m:s]ù��K��)����zzzU[�?GG��#Nwu"�,G�{6�O�{�� T�j9|������y>�ϔO�&�!�o榇�7��E�(5 ��Yvw��@���I��;_58vb�]F^�l\F��2��Y���@��d[�{�'3��i�un���M׎�r(�֬�w2N�^U�=�n0ڦ&3-������1KGҟݹ�.��N��1���/�2c����=b�o�S.�|pa _U�����J���՛͵}��]S�g�|7ȏ��7���1�T�������m��ӯ_n^�����x����5����ޣ<~��7��칺ۿ�>��m��u�����ډ��7�1�d掫g<2`�KI.�U�y�z�T֫����`�?������;���ƪPBS���	.X���5��$��5G�fƭ,����@���0�i��h��T��ȕ�b�j���p{�2ngLy�1G q��	�^�P}�|f���J�:�j��qX������*R�Y�K	��r�[R�<>���"M��a�O\��Q/'/�R�����Kq'e�4>s ]D���-���3119�X�W��37��l�rX\⋀����ܞ�KߩJ�蕭4s&UHz�]AR"�/l�`ط������çR=.c�ymmm����i]c��M��珛�9��wq�=�p�%%�B��8�<��2O�� h��]�`.�<P^��,�ţ�W���H�ұϴ�l=�]�a{��S���sx!���IZ�7(����������#/CKf���K��-�k�~(��8{A�H|]Q>�:�RTCV���Xq�,O]511������̲�������.�Wn�	Q��v��G���h$�\F�h�=ijj�z`�|W]]=U�fz�>6���W�!\ⓣ�OAN���bf||jT79���-�C�d ������]7��Iu+����:�vX�"��>�B�����1�)�h�����|�ΝS@l��Ċ�G���i@�������mQ��Tju#��4x���P4�4�:�K=��0mV���u����M�z��?Hdk���l-�,��eKe1K��ҁ߫l�Z���� UD<�&lߍ`L��,u -Ҍq�Q����	�TaS��ȫJ��=�?�_�,��f�����a�dWkv�ڎ�A���ч t'n�9ȜR^i>z��(�Y!uԀ�n�$�`mr�J��gl����I�X��f �}��H¤|�p�����^\��g�K���!��k�/�\��L���Xb�_2 ���]ȨϽ�̴9���@}�w��M.133�;!6XX��C��Dk5L�!�ԯ3H.G.��l[2�/�2p5��D��U�VەURV.�,B���1����'O�e_����L���Z7ZG8��p[饐�����Z���t�lF���O/W��0S��v|!.S�1���E�!L�d��Ɏ�<Wh��kk�����w`;'���K�Ye`�?��D&f�e�	.��Q��@w�/1���,OE�W�JW�!�-g'O�<U?����;]f�K"��CH�uׅ��h}�=i��l����V��.�x�[8��۽��e�.�D������%��� ����}Z�-���2�4�B����|��j�`�Օߕ��g���>|h83�Q�2����ٰ��v���꧹��jr=��J0��R�l�������/--=���6y�|�JfVV����r����W�x��Ek!�����?EN>�ʞY�fe������}�V��d��7]�tؤ�G�N�ɠ�N�?���2�nI��ޣ>S�dd|=�pu�z�����5���}���O�uu�jjj:���,��vU��E�$����'������#�$�������x{jû|��o���f+�p��:���,5�����s�MA,"��w��_�}w�����d	�S��}�w.�=���l�H�Z&"�����d�~���}������%�:y�B���~0�y��(tL\�qZ^Y�x8"�E�!�~��,�(Y�o�cn:	u՗��Td�nmI,���57�����9{x���Q������EB����˟�����(8[�[��A�豱��|�)�� V�����AEN���,?���O ����=�8�&�4�ɞ~�:8���qΊ��cà��i��[���,xg.��x)n�����%�}ڵֵ<u�r�;�WJ��`��l�Z*��"�$�����3S�΂�#�F����̬ �־~\�JKf�k�w�����p��p=?Ԅ�#���O�Q�M)��h���#��"�=׈~�N�|������V��d�lg����*���ٿ�f�_�;�Lm���v���A<	�����uz(�M�W��$�T��o�o����#�55q{p�Ş�k���ZG�@%����!��,w� �
��� ��a]����H����)���T^{,2���������m6.����l���#�SZ�M��0?;������۽8�=i	��"ps;���g;:R�����!԰( �W緁�1��oTH����Q?�|V[�x�ؾ�C�;���CEM�GA���3G�>���CD���ڹ��ǚ��1�"�����U$���we0�+!�ّ��HnTG����O�\�u����]��;�����Ilf/���@T���_rAt*�d�X7u�8�P�1{�r"���҃|�+k��l��\���EMd1��C���������ײ�rt<:�TwZ��B΄�Uq�IڠL窈��(�t)�:/Z�j�pJ9��j��ׂ�¬������K��b5��VxE'#r����84�5���]�L��Q���4Il�p9󅊓Y��T9��w�����t�)�#m��;�;<&�L%|xH�����Cv&)I�mv�gjXa7]��1=��#�l�±o7� �sX��&M���C�ޑx��c��WY��5�ޏR�7m%id��
�!�_kVA�4׉��,��]�u�R�@{�I���x����8,lI~9z��^]qp�$�ͣ���78o�����d����g��Pj�
�K�D�}pg� ��X�"�lr�"_Ѣm�韴T#d��KA/fI�.�|6&Ue�r��%.�T�Ti s�C!���w��t�>�x� ^f��
XK����.'��ܢN��Ng����%��r��n��G����O�U�u��Ύ���e��|�JUg���gz�:����l@����ظx4�:�u��%yB�!.�R��J��T���
�%p�w���e  �i��(Պ�CS$������U�Wu(jn�oܨB�5����Г#�	+�k�������P��wo�(��)��d�jW�x�?�[�6���=cZ
!���F8}��H�=���TO�'$2�z���*����?�VA��@h�C���c@�{oRܝL�۲[�<L��[�譊��E �VL��Up͡� ���d�RS��*#�>@�o"8�t_��1���_�wxr{�@���GY-E�N`j9����N�|��_����Bk���A$t|�j���v���W"�2N��sﭏ��{l��|Drܛ7oznL6�~��:p݌�����A���^J=�;w����+*&�z��f܇���i�����QI�r=(�3�#}Mxؕ���$eh��(����fQ�,��%�ث.�Ш�,��=~�AW���B!�{Y��)k6_<Α��[�ML<�oʿ��ɓ<����	c��>k��m"�KLL�M9H�1��r��P��/X��?2��mq��_�/T0���������WS��i�Ke)_T�X�� o{�.�"�>�Uz�T�U��x��i������#|�N�<���w��{w���8���e�b��pA�.3[���h�����j�k�F14F	 �4;+�<�ya�cV|�%�$N�!Hq�լ>r1��#G�J@ȵﮡ�w��l"B%��^��W*��P�z1Dqt�>F�[����/pT�_���n]B^ N��1!�T	�1R5bbD~-�ލ��j���Ji�Ԟ���C��KX7��"��<�[$���XZ����z�����ݽ�x���vu}*����h,�u����+b���aϸH�i��A;�|R@AO����z��|��O.�ǀ���
��N���N*8�/�����ܔ��}�/�؏�y�n�E.[v�M:,�&���`k�m�k��K���T8�'W����62q�Բ���tB��]���^��>��I�(HT{i�aib����Kc'�Ͻ����j��c��i�<��A���ҷ���ڌ�_�``�_+̻�d.^�1n;� �m��q����TC�,�k&,"��u�������ǒ�`j�5L���[�$ p�^�,Q��
�b�{�F7:ÄVG�_�ɴe0����x���d.��]W�f�#�2��;���,�$.'����@g;�q-��cء��2yڕ���#KgR7�����&�)�%u/���(S�{Lv����l.��y"��T�o���8�x���MpPA29Q��M��>K�����'��u���O	�K@��
}�;~V.�*@>���G����u�'bY��zC��.϶"�(��+M���B{"w^��V�A���KR��)\�ŉ�w�s>��+�.�n|�nBE��'5ϸ�D���8d��a(��IC�|5@��:G���C��.�O䟬�	=1b�Z�0��' �B��s�wԧ�{�����"#����%���qe�q d_4���g��m ���׏��޲R	�)C1�1_��f���r:;;z����U��%>?��zL�bD��h���bMLLd[���3��;�P{���8��<}�����R� \��`���c2�:��?�4�"ʽ�Bt������u_�3���w��ܛ����xo�*��m�WI`�����ﾸ����W?��X�Y(Y���e@/��yo��S�����vޤ�� ���8�q2��-��=����t篡;ھ.G2��u�o�'�>qr.����k�	ۚ�e�ݵK�s�6yް����%�� }E��ؚ�se)Q��~Y��<ʟ/��/o����5^C?�����E��~sc\�=�dt���5��}-p[������(���]�d��A��<,���W}��xh��q�4��]�aF�y�<�|�"�́!�c?����1	�ac���MGfq$�7
D���-�,�W���jk_!Z�a��p��}�˓=;d��W3N�����9����v{Y!3ߢȸp(�:<��\�|�ߺ�"i�&?�zo����z�i3�WXޤ��U�:��-gj27	�s��
5N���ͺuX���ҲM��r-��
BRv��Vʉl,�6��&�����>�У+��̼?ނ&�`#>�؟���||���x�ΐK�U�6��ߨ���T��U�y�m����郘E�&b��3�����qi�e�������_�s�c�>5���>�x�G�i���|AҒ*ш�}�M���ܣ��YA�*�9z�h$��
6�QO��P�s�=xF;�)�ؽ��D�5�{��������P�ˠk��P�;RO��b��=��[���Y|@*+��?�AG��ׇ� '26b��S�znF������A��:MC�ȗ��2'���9���J�繋��1�.aKo�^;Gڋ���șF71ӑ&���'$���W���|�����h�7�coM(�p�[��H��W	=���i�g}�C��D�O�������v�'e���s�jTLw�ܴ�<+�G�E�1,�A^�=O�߂�^"�MV�?�7�&��.Ad \���/�$��Q�eD�s��&s�#8;�0!�V嗫b�e��p��Sz�ެ���)��L�ʋ���wz�=�T������U1�6w{y�]Z���d�n��D��g�r0{����?k�q��ۄW��Y~ N����О�Xu�n��i��	oIy��r�.����/�^<=~��+A�J�_�	�����{�G0�'����۴j\��3��6O�$����& ��Z�7p�,����1��2���9�Jq�7*[���� uѷ	s�R�|D����M�1O~t� ��<� M/�w�+�&=�!�ܽ�|5�7��J�a~�������\���<�p����m�,������fy�ٗ��$k�h���D�[����4��������$C<�UO����m@�u���u}t�<�e�����"�Z	7~xm/0S��c�@��&܍�B�<���%�.�p�?����"�A7�9��m�:ٹl����C���te�4hkA�����2�jw�����)�f�����ku����&�l0� d{�����se�wy(�����m6�v.��.��l3��v<FkN4==�>���� ��9셍���b��h�n��/���q--�|�r�D�â��z�D�q5�0c�d��/�<�K�*���ᴩ4�8�"���@XcA�<p�3C���0��3iqx�IsE�g�A�#�ר���(�i���S��������g���I�1��m��A�_�`�klJ�㦌K�l��70�Y�h1�X2���^ƬX]��=�5d$3j�0c���hӿ��ၽ=�"�C��C�h�h�	Ԭ:���嘣KKKe���g�O#l�.�����SR0 0��g�Я�l��LRg��(yˮcH����,F��i���Z�q��;d�b����<����n���s�ܡ&PP�8�F=��k��o��p2{��]�E]��	�����G7 (1��{i6���_:X�'��䙥�u/�#x`��z�߇o��W������~�;�Rjz|�ֲJR���((-YS�e� b�]�*��/�Ik�n��j8����^���14:Q룜�� ���Ǫ�N���������b,]�1,��#����yӊ5�}_���U���3�K��?S�j	���Ls:"�y�0 nk�E��܂��X�T� o���P�7��p�a�T�SN��N��=�>�Vf4|4a�����L���&��J�86��%�8�)�I���-���y���<��֤�i�0�Y��@��^����u���2��8�<��x��)�rD���e��.�`t���\�$ڏ��T[8�^������7�V3첽������ruNZ:����CM���[�[���cEi&h�"�wê����R�@��uh1�a���7��\p��묢�;&<����G[�W���9ý�u�����d|!]��i꺹r��YGiN��^.�������[,���|<�ɵ���e)��V>��u�v��_��W�GQ�3E���r�
���d9����m�N��n�z����z48v!�}Te�pB���D��=�z2{'P�*R0����B�.JݺAUa�3?�V��
������DP�[��^g��X:�ΰĢ�Mzu�/��ͳ�G߅Xb�V-�UC8Ƥ�#eoOSqkR�1˻��X�?������5���<4�l���v�4��b�'� tvnn��RȜ*�7;܇Q]��~� �b����䛰5;�
�����x~��l$t�T���$��5��坖uI���@'Q:����l�ʴv�_�ت�.0�f�j�@^�o�m�.$<}��%��y�Ȩi�T&!���-�J@սT�D���I
�FL�T7+��'�-ɽoU��F�樨G$ O))�=��~/$Z1hM`������D��P�����2����4���;p�[��{�g����A>1�=i��ۉ7�iFL9�C!���̞Yj�P�5e��L�F�������-���Pn�Nx�GL0���}��5L+mn����x|íb��;K�D2�Ġ�p������F_�Ah��'w_�����Z�T;�������,�8X�,�>p�iY���7n�i�/7??@�t�a*!�P!5�p�׼Bs��?��s�jNf�ϕ�� ��Ƈ�9��X�� L0�J�6�F�����rmu׉g~��"�7R(���nhDۑ/g���dH�@�)#H�;���k݉��_U(����n��'M]��a����]^��'_��R�M��#������]t}��aC�hzz c?
�_�wXH^�.�ዂ_�9��D.l�J@>�/�}ت�V�4L�U�=j3$��&T��,t�ѹ�o���[9֝.��/w�U;�v��s�b=8[�♜7��Q?V	��W�U�Y�ZP�x|��������������?��q�����>��Nc9q����sݜj����IU󳊆�D��	�]eQ6�,x��6fLc�j4�/i |>ln���D�aؒ�l�����J��1a�Tˀ�����Y�*Θ�ʾ��m�^Jhh���H�詈�d�j��O�����R��K��g"h���s;�i0}��u���>z�W�*�H�Ɲ'����h�s�o?����^��@*�%�E�{_��mddem}�&�o���4���YW_*�<iP�v�+���o�"Eg�)E���M����KY�=��?��R&�4"}d{�����7��V��c���(��K�������l2���d'g\* ���)mU�Z ~�����VA����;�Ʌ;3#��
�s��&�����\t� �q��Ș-PX�|���ѝ"��ՙ5�ض��ԟ��%N�뜞|� �u�x���D�d�����Go������	�������{�����5*bz8�eb���R"�0ziQu�����0�Q��b��H�͓�������.��k]u��ǝu�KW���]f~����Έa��tI�fq�'��/+����&����q�44�׳z' ��mUf����0W���!�z[
�H̙��.w��d\���#�>���JJO��xlO���Z\��cߞL𤐽{����W����f���(^ߚ�<��vH-/+���$��n���[�la{�o��{���%r�OY�?�v|�F�?I{�B�;~ ���[ѭ�q��&�4�o��YjF���g��S�r���Z�$��P�2�Շ8Xji��1IvĿ��67Q�t��ͻ6���͓D����V��ǭ;��E4�S.ww�i��?,�Xv�V�*0em���uu�'��}��*� E��!Y�N$X�#+:�=�F0D�K@r�I�Qr�#���pw|K@�Ge�����x�����(!��E�M�3D*#YWF��q�k${��ɾ�.�ȺHH��^��6���5��V����xxؗ�=�s��u��uYm��A�|jt����D~��ƛ����ƃ�\~�'�|JP5��6s�����7��Z�/ �d��]8���9!H����i�'����)ke���	N��y�_r�&�6�֭�mD��zд���=P���\�ᾱ���ǈ�P�ڥ'a��ͭ�`D�_�4#7g<�i��?`-��}a5��>�YO@7����<\���3lMm��`��S���*��IZ�6��8����W��ԉ�l?�	�^g�Ҫ�V�����H�ݙ��sÅZ𑉷1�S�
6���}<����O���R9����FJX;��L����bV��ٚ:�/xM�������M�|t"{���gb&S���te�Ѯ�P��������	B��,a%���<��)Hp@���~<���u�����NR$g���n :��4���bT햹�2�+5�'��~/�d��~��E��
ka�Z">�[����3z)��:ŪkgG�Q�-<�J^]ݽ0*��,��w�����q?b������}ݣ�[�nǾ݆i
j�J��+�%7ا�����Qv0�~~��+Z$j�p,����H�}�zs ���p��f�K����޽E���cF�{"���?�>�\�?C��5�X'�%Fl*���7>|�A�*��ھ�G���������O����Y�:N�i��;o�4�F;@IJ��򒪊	��s�
��	��z����y������״�e��h���f��FFc�N_���fV�~l�me'<���Q�qs�JE�༎x�[ )�1,����ZgbW;U^�1V�Q��H��8�S%�i*|�'�����eC�G�P�p�5�?��Tz��-:6L�UT�;	S�;�۱��)���=�D@�ږ�`���n�-����ȁ-8�:�܋u���~U{s�k�����NA����V'\�U�w�uL%�yLF+ϋg!"q���7�Ŀ�0E��U��uߴ�}��염���vOZ\@o���~�ư6����r9�HzT���k��9����D�I�N�34��-���8��N��NDT���HT9@��&�+ۋ�̧|���Z�H`ܓ�#���-���x
-�b��D�I`�6��{�B	�K����I�3�����^`)-8t����6(�E%�29y�OD������U5�~*RI�RG�	�w�6�$=�&2x�pKp�ޙ�24r8eLz��5�U3Myp�x���x�g�������F�B`�Sr��Iu=�fE�ӗ�I�'�����>���� ��9IK�g��y��6̜b<ot14xϘ��C�[ �Jbr[j`���S9�ן8\�aY�Nֿ�;j���[ ��=�\,�>kx'QtZ������|�;�u�
�R;~�Xo�[����K�"p��b8KMH<���)�K�����|����%���+�Gx.�&�����������zߑ�D�n��`0;���{э�?���F�TLY�_׈�v���>`y�W�������N��:3��/D�7U�_�n[b��zj�RA�g�F�����~���]�)�ϵ��*	l�da~an��7�hTy��^�g6����2xn˸
'im�����a'i���3g�e���`��͖U����$�((ɠ�r��S���U	.ٯA�b�6g����/8�9|���ǫ��n�%�7��9s;�u����V5cj�~��$��R�3B�V8���{�éhu������c�掤O�=��~��o]&�p�'�:H�{�ǡCM�IF?�0u�>]�����47�mG[ݎ��^k�>�UJ�������+ˋ�mǢ��z��q����oC�����v���jfEܽ�+�=���|�у��^��_#z��ܚl�Q��Ͽ���x
9^��� �^����V��gNI	w��ಌ�3�NDssW������2(k��� �i}���_�sC0r���y��� �d��~�5*���1i~�+u0������ s�ݴ=1��u]�z_�OD�s�Q0�y��n����ln��e܊�t���zI�#�~�$�k�g>�� t��ڂ�P9�J~�́Ć�h�2��lFcS������&��c[��.�G�Y��z⹀�Ŏ;�k ���o.�� �l�-�(��d�Q�y�ȕ���7Y�1;�:+&���k�"�V���z{�T�hJ��,{Ȓ�F��1i�,I��Z�~����0tmn��H�T�QϠ�2������e^�m}��V�B3�#�r�1$i�ۡ�=C,!Α���ځ��p���7���ƛT�S0�XS�����*} "���f1j����=@zA��p�P�������:�ܼ6����}VW�ɲR�S�u8r�7/f
���M�	Y�Z�B�ùT۸�C�~�%�Uܙ
���ݾV�v*�l\��G���?U_n����pV�]�LW��y�p�6�y�3��TGֳغ�������}V'�b�=������ ے^��vV���q���F�9\=]��Ǜ���:��*�m!턶u�m`\x�^�s�J��k
}Ѵ�Vɹ����>Ҹe>fW�t/��6`��^U77+�z�DMMmKH� Q���)�n��2m/_;�?��Ư�hٴ�zr���f���嚪��6fe�c	������c9}�O���d������	��P�1�B�U��Л9�Vg�����*  ��K�k�����BTTT_p�'�+�R���+~���+�>�Z���~�*..�/۱��m��-,�L�"��z
�D�5ɪ�h5 _q�+//?�����N�ş��̍gc,�认��CwQrq�q��Q���)�t[��)nf����f2���3^��m��UNp*|�^?��qb�CÛ5g��.���i�c��"~ Bt\��B�I�Ґ��V�_��u�֚j���Ό6�)�W��Ln%j�/%DEC�v��n�͐F���$�.����}sf\b����
3�9�[R���5A����$���GMVI�N���-+�B
�S8y'NNI��z�
<�p�����-���?�N��S9�v��uf�D�;lλ�o5�7�R=~5��
?gH-�8BM�qs�Ip�-����v��Ru�Q���cdB�A os��5]��ocI^7�Zgٞ��V�=��S��:����˛�Ξ�}��+����2$�#�gK�m�~��U��2�J��GU�0��:�����J]����M�2�<��؄�G)���Š��3ζ���BWשX���l�m�=�2=$�K��������@?�V?�m��~Rv�{'B'm�9؜i�!sn�@0U8p�dacc#�B�É*�����l̧	�}����������ߗX6�
�^�����1�R����#�W�9���`��Q��>�=#*��X�c>�x�����b+��E�+�<�:�<0���@;�ug�*��싞�����l�:\[��h�8�d��v�K7t�<\�A>��i6d��q��$]Ӻ�s������J*ԋ���ܹ��d�=]���.�jv,��%]sY����C������q��B�l	���sQ�K�9ʹ%.<u��������Qr��4)B�v��=���n+{��&��2��7m�L�m�3b�ʶń"�E������Sљ��AZZ����z�ӊ����DYTLlع��׌��羅������!c�Y��������jDsHp�:a|����8�������RX��y��́�'Y��Y#'�"?��͔��4�*��x��6݆�I���RYYy���8�tB�����M��v5rI�4��yi��7�_f,y_�/<}Qy�
շ��j�`�׈�/�{��s��9R&{�g]��t)�W&�ʎ
U<@tF�Z�o�4e�!�����nK ��e*_���8�(#���*N<_5S�����g��|����X����G���r��*!^n~O��/�iw���T�'���2�e�pu�fU8��7c�Z��S���=�O��!	��E�S~e �j�͎�OZ�w*���vǣY�=�Y��	Wם��f����IZ�1K�A۪���;�n���Dz���e��ñ[��c����Ӻ� ֺ���S���ӷs�(�3���*߾�da�]�m|�,U����CzfNM�hN���=$�8�{��rȵ��u?�s�z�����B�rӕ��H{�y�VPљ�洵�32�!FGS[  ��H9Q����	ݙ�i����g9��������@v�l�����J�v{�\f��k�.����,,���ݲK��6��8OЁJR�*����2���b;+ߥ���u���=G�Éҕ��m�����RY	��fj��G�~n�z�:��DY	�@g�T�b������[	㑟�nm�\�8|��ƙ��On�Vf��x�d�c�v�oL�b�J�S� )=n�R<e����.η����1�k�34:��m�;���S�vf������#+���e&)�E���ǲΩ[���0�z4���	|��^�_/=i^1�Xvd��c{=����|���l����腶S���ں�Ku�����N��>uW N]%c���7�6��/IS,�.'-��Â'�� �k��1pI�6UG����vO	
���J}�5��_w꽿�� �6/��;e�5�8��ƿ�K2��"��XU��e]8�:Q�xM��'����jZ�jh��j�&D��K���S���G�SAx+� �kڔ�����c8��õ� ��yk\+�[�(�3����N/g�7����%ܖ%c�Wm'�w)�%�g�Bv0����P)W2�nc��Ґ�]wrDFޓD��҃R�h,�C��g���:��O������i��B�,g�be�ј�ũ��6.3T���׉ �M�%�_����<��+��qJ��zR���y�'?�G���E9~��բ��U�cK����������Z)�=I�p*�EX��P�cojaV��M�*�#cD��&"2퍹?M��Vt�aʭ���4�o=����Խ<��C��&s�Ȣ�5�����j�p*����/�b����g�#Rq։���$o�����6���Z $O�S��:�hy_%%�� �~�B	���XP����Tu�v��V<����LIu�]�e�{k�����;��Z�	������1��R��|x���3_I�1���[j^����6����8�*���-���_�2t��[��z���o�@8g�ž��C�8�RܪSe��RK�r��M�S\���qK4��������MJ=�T�+v|�Mj=�b��~#����� ���Wn��hH�H�ib�B0�G>�ͩ�,1v�����b/���߹������J��/$��S��Ho#�7���ܵ��_(�e1P�c_z���+CZ�m�(SO!�lz�rЮ���d ����<����_�`J���N�0/O/}�T�Dv�h4�;z�>�a�"�\/H����jk�}I�w��Χ) ��v��{�6��4�Ѿ��Ѷ-&U�٭-q��tBv&\��b��Bi=�P��5x�[�F�	Ug�<o|z�b&�9��C�Y��G�q�n�|� 7���6]�El�סw�c�r�ǯ -�L��9q�;Y��۝�;<�}���6���Tn��f�M�)E��1�7
��tk6���:�Qɷ ���^�w�#�*����Wk��qK� C��9L�I�=齾��W��s��(~��ĩ���>�zrL�[V �e�㥒t�	N�gcN k���R�#��Eס\L�R���A�����fkv��\%��3>�8�KwbA�Q{���}���_n~~1�cRP�A$�.��Ս�RbЉ�:&�e�\�\�o�x�X��>���K�JH�!�}��Dj��+��������+�6ޝ�{g�s5&N��s�0cf(���hI��0�v�P��]!����I��U��N�vtU+*��P�R}�W9~7 ���XΤ9Tp=!���*Z�/���:����E��U��k3q������6^=�'Rʥ����iQ��<��f�V[�WZ�N���y<��p�:�u5��s��,wy!�f�Yb(H�!o��"͐]��r.q(W�M���5u��D�;�����ۻ���r.�n:Av/�ĺ�,Y�*-����I?9����m�J/�Gu��+VRm���=Hs�R����S���t�u��U�?��^�af��J�c{��:��8	TC{��C��u���#q�Y�'���g����E�~��_�SsM���C�iB�v��2�$�c	�����V�/<���`f��[��E�l�^�����d��H1�Q��aN��-F�X�hoE:�\�Zw��wc���6���'��ϧsm碃<��'�o�GM>J�>�#c�;�����c��DRH��/~����T.���%���M�v@�R�.O�Ӓ�`��cn����'M�S��ͧxm?f�F���/
�*�=�-ڂ��z�@ϩ$x�O������k��0_��z�����x8Ŝ���z;��R��� ��/;�@s��F^d�2;��:=���ykn�@.F�r �Sٚ����,mx�C7o���әtz�t9dc�%�3&�����)u��|����.�@����ka�#���^��s+�B�mc}�54�.��/7�r*�9܎�Y@��<	J����[7��pt���Euk�=6�:�%���������R��8OC#FP|���vqc�y�?!O�ڪ�@mԭm;#��*�E`��oOW����Rd\�./;�y>���zE��)�{<	�X�"-��n�"M��5�#�@��R5ᠩ�	�[X�&�3�Q�����H��"�Ӓ�I�j���M��~���%d� ����Y�(������ ��>��;Y@��lY���C���g�s{���Ar��H��c���Q�l4r
� �D$��}�]K�yʺI���m|��o��g�����S�������߁R�.��{�rP�]������~�y�������4�ב ��ڊ�l�4َQ�i��P�q�Mx��T��QJ�淇�zƱ��yV�
*W��'�Ķ�p�xy�mf�So��x[�l��������ކP�6�!�-�þ�P�AIP�� ���~�����!#M�џ�T�d�T�T��|�뎫��8%ů<��/��%�F̪�[��f����禔M�X�>�z5j����׍�v?[�����p��}Mp�U��F	��,S����m�Ej;�-G��n����������pD#����o�� |t��]X�D2޴]ІK�����O�4G΅�S���~�H�����+S�føĠ���:�緅d:�$�|�8���H���p"����3ox���%�<�s���Rc�ܞ�Q֯�boq�*�Og@��UM�F��i� ܪ��[��xe���	oW�W��s��x�EF�P���f�	�G�q� ���a�{��&�kc������=���XF��B�>�i�e��?�$?5�S���ތP՞���v��]dN�_l'�^p��c�=Z��\�+�;�6�'A b[Ĵ�,%��3e��+��&����)��؅Y� l���i�>�*#t�@>`�,�ʏs��s����֖�ɍ7^��١��z�F��~ϧ�M1G�!xY����G�D��RrZ0�p؝��KO�ޟ��h�
�.�*��@,ö1��Դs6;tW<@&,W��deeϑ�O�<���B���3\+���Ԟȁ���PQ�$ơ\�
1����"������������[�w� ��_��m6�:W~pW����� >���$�Q���$÷��ͳ���?�`�b�l�ܥ��3�Nnr�-�pt�옐����>��=
���J(�`�"ں�ܶ��v�^�_d*>����)H)���\�||�>?| ��%W��~t*����B�s��N�.��[$�Nﶟ��F{��B=�60�Q����[h�`n�AR=����@KN��	�o�5	���i�PF����S73���G	h����w�{?�zw�$;��������|^6��~g��O��b�o��NP3.$�>U~�i�ݵ@C_���j�
�,��7��y�pр�6���=�����s.4�N�_�]��2ͷF�I7�x��� ���2�M�vK��L$���u�Y��:`7l2��tMw�@�I��\2��}�+S~��N
���ag��y��r�*���tSs�����| �Z��լ��
$�8Ri����n�Cz�6�]�	��/Qg�+gH�mED ���!�5��Ԛ�LĤ5��
q���EJ���%^��	���m !��#����R.!{t�����5�[����j�@Y��K=c0^v�b_@^�_rmOY2�^��8M���g+kT�r���Dt4s$�6d��ں�T���:g��Rca�t7"��yxxL'_�(;���d>t�؞�!3�$�N����Ǟ�x>;�U��o�u`� ���)�L��ǜ>��D�u�W,X�SK7�Q��^6Z���q�j7�9=�)���� N��kϭ�ў2�@�qժ�I)�PSξd4�<���q<����������F?J��p6�PeM��v.3�D����Et�L�;�D-y��9���wd�)���@�+؟�T�{�|�u���[|+j`�oX�Qc��M�Ҙ!p�=����*ǻ	vN����1��?���G��n�neZ� a=�s�â��ׯ�Q."����&j�խ�VNʒq�t����r{���G���O��BE �[���4��k��T�j���௘O��
�;i�'�g�w)ֶ��k"�z+�}}�v�Tk��=������v(����� ���p���*z��z���K� RaB'�5�N��]�\�yr���S�?��$y&�4��v߂�d�Tn���S	�����c��7p�����7�ꅅ1����C��{xߤY-(S���d���O#��J,I���צ���|mƙ���$�Drܙ��������'r�b���t1s�k}�'���F�񌇋�68��
�������.�J7�xQ8����ܳ�F��1Vy�H�߯;z���w8h�Q&9M6�<�]�F����k,�-\��@�A����fk9� z_u"��a�wW��JH��)7Ag���V?I({�������{c]{�n 4�*�l5zZD������%A����Ĭ����Ҏx[@���$� ~I6_���V���d�������߼�ww�$�}:K��4-Ѐ�{s^K����L5��6gv��\(w||X$�}� � �z�OD��GN�я���j����{�#傋}C$T#
��\��aY���g�d�ͥ�)�1����NOt���4���lڻx��vi1�=��HEx������IԖ��؈��cf�70�Q<\hO9�ٻ�c�+�̳��6��N�Ɩ]��<���f!�1�"��/�aPcDo� �j.����e���D�\U���JD����E�\`yH9�L��KA?�NO��C˳��=�u7����ڻa�'��a���m�vª -_���C�\��p�l��}=��g���f���4K�����X2;&�Ű>��6�;�ձ��r�-���{�dP��v�b��SN����ꗟ���Y~�<��9"�0�\���>\���w��;[����S(��fw�r��Y<�,�PUJ~� dS��5�1��G��~|愞��>���o�io`8E�L��;�'�k~�w�=���D(q��K�6?B�׿�Zn��L֦����H�v�U���~���!��;��MB�����L�Н����_����IX�e��e�EuSk�W5�X�s$zt�J�Cl͊���4�e1�?�*���:�+����,�P�a��Y�؀���F���oT<�[�ne_s\���/�,��K�җ����Ir�i�}���^�����O �i�.(Oz�1!�g��>;�o�(-d�l�c����#�A�Q#�����ZO�*�	A�$R��]��l=��&)Ӄ?�4��2/}J���{� ����a��ۼ����i�%D��@�,�t��V#�(a����F�%Եf�)�l
�ߺ��@%{";���N  ��h����(\�
� X�]�ͯ��a�陰��&�!�2�D��x�k�9�5x�^<p�_�]c}f�<�P?�t��a�M���W���o�9�t>�-s��\ S�sw�~YD�	�g�B����)Zm�b�@�2&�X���)�i��w�P���<7�G��̚�۹����7S�k�ͯI
�@d�B���9V�Ց��q�e���2%1VY���c�M��1ͷǚ�7�v�c�+Y(�27�/�����!tA��o��l��짲����'�ާS�lz���X�g�(�=Q�;Q$%�w�e=�i��C��
3�jF�~��0VZm��.�)����ذ�5�ʮ$��,��V��0��JeX�"�u�!-�cV��M��:�����CgV,��ge>�<��i��ߠ=�BG���&��ty��f�xG����̐����I,X��㪛j������H��'��ǥ�>n (�0c(��f���9r�����7Dܖ]�$<-T�q�.D�rT
��opE�l)�(p���m���OW�޹��5��u�<��b��, �����G'ʏ����	:(��<�#�؅�<�	�:�?z�m�>�H���-{�E���e��t�ڟj6Dt�O�\<%�:�������{��������k˳��c�X�vln[`u�6&�Fb�HAI��Xl�ae��s�;����^�h��o������g
o��x��f���АJ�{�%�_����� �?�`ػ�$�[RI`k2֦M���`���gxO��
Z�ez迋����
)-��c���V� �_�g��rœt����hrU��3�pM��徘�~~�U!2*�Aj���H�7>|Si�|Ǹgc�0HI���!�}���OT���Ӳ�t��k:�t*��S�U��ƫr_į_ˮnr������F����n�r��Y�}/|�υtGM(]�?�[���R��SO<j(%b#,�@t!xR�-���Y��'!�7�	�����e���,'��A>yش���6Gb�&)�����{��7wí��[�-�tm����'��j��mU)��e�U�1߸.�"� K��C�z�[����s�'�l��;���}3�)�v�"��,:���Y-j��7@��k�����z�!| իL�KE����,�;�\ɵ@fD� t���VhS��=��i?}}r���:����Dc���%�'�Ye�s%)|K˵�y�iِ��	)'y`��V(Ab����
�"In6vp��,��eRe)�-�I}��'aJ�߿����?�!Ȳ��mS�'�'����~��ڕ"��)�u���yI��q�*fa#wC;e��w�V^NW�.�ɩ
Q;���
k��I'�W��
W���7��D�1��H�Ԍ-^�^l*�>d�*���{JU�@��ڒ����@0%$�İݣ7���ӭf6�����ί逪pt���8��:�-���՟��,�Kܳ�o�sJ{���x��5��GL��h�W*mF)�P r'>G�<�<b�3���v�(�5Ta8��;D�@��6�u�/$�Ig����|��e8�qh�i��Z�M�R4�ip� u�tak�;��Z�i��a�UwFk�&X�b7���I"�Eg�Dq��?}���C�a$�CfeS���v�ҽ��R��w4���������ml�Z�����[�A}�cɝG0����X���_)d������&�(��/�&I���u���<���^ڢ�{7���ZsA�l�]0%���h�8�s�P��X'�m�^�-����Wў�Ȇ͹�B-��A��1;6g��@��%l�d�׀z�@��fX�x��vl�K���,O"r'j�H�����<�~5��pl��S +ſ����w�V���4[ �fe�Ti�}tC1D9���)G������;�e��E�����l�{���L��Ћ��|��50��X�u��]I��K���b�\���_��
�7z��n��;�j,R�����<&C_OA[�I<��A��"MnC��0_�⤻�و�ޮAZ=��$%�N����19���ؓ	�ՋwW1�����UH�V�I��m��r\X_uI(��?����+)��*�d�壙�$!.zNذ����N=�ǫh�V��ϷR�������k@���!�jG��K* ���u�߾�$AX��K����f��ϔq�B/�p�ёE������WdK������	^`-8:���xl��K����*��ɔ'8�:!�������7�!_�v���v�'=���F���<w-;F�p.Et����[�����L-�%�''���7Ypv/�'VU6&���wR�!�)M�7��Y/��r��Z�V�\�_�~��?��q�?���(s�sn`|�$��6U�JX�z�H"7e�_�б��5�e��Ӛ�D��;	����]s���G���!�a�P�������f߂%�j|6�j�^p��%��R5�S�b����h9�j}����Ȑ����p��(g�Ō���̼�ю�g���E�ƶ���<�&͆���һq`4q�Mf��,yBt�a��+m�ڶ@�cў�i�iX�h�$�v�3G?���<A����e���'�Z�Z����F�ō��g��`f�s?
��]�� |�6��x�]��a�ҟ�����}���z����I=ˬ �չa��Y��D��*t'L�?>�棎���=I���	N_\~ݘ����v4�eSoHqDZ���y�z���PDU���5t{��>H�\*1����z�	�*"_�����L�!�����>��~��eô�pȦn\�֎)������,5�R����}�>��kI��kt�BV�ɫ9���1�;���@gvh@\�=��(��~��I���rOOʿ�����կ���߿��]�6����C��mY����������5�d&�X1ӄ�'����⥵����ݏϤ�[HNu��ѫu�!�����M�*���"�Fv&��������8><�/5�-l�[�m�x��c���!�g=0  (�*<��X�0`�(%�����(��r��w�xq����|�v�<o�J{�;�A:�/�ܧX�����Tf�1�����U-�� ɛ'ɋ4ck��q���������,�L���Uz�u�PVN�k�<���/+:D��ߦc�Ñ��Z��lO�4�`w++(�rzY@@ to��
Ao�<��%����>
إi�3WK�'�O`���I'���5�a�n��̥�I���7�ă���ݝM���i��+����SЩ�9��ϰS1֥�_����3Ks�*,��e��h�Kk�6'88�� �e�`���NVz�=f��������G����<���?u5�	���,,T�;�N���{U�R67�����6��A )�E��ޘ?�J$E�nZ?)C�e��8�&3�U��E
/��Kr��K��S�U�Kz3�Gi��o������&�/E8<=�b��:8O崹q�UW��`�o���}q�'ؙ+3�����M���ރ��߸ͭ��S�S���~��u.��.�R��k��H�)�륚��G��T��lݘn��[��<��l��+�*��3���=ϸ���g�O�GVH�6�9���C���`���?�p��x�rJh�|���S�h�aW~��.X�)4!���7���1�=�7��c�mG+xe�lڍ��伴gnE�K)�[��rV+�#x���T�\��'m��ڜ<ɕ���ѱ��X��Pӭ��Ŕ{9��H-+����5�m�ޖ��/}�Qqϒ9ޚU_���t̃WOZ���$C�g�_����ض�)�X+��(~� ʃ���)P�?r�$��_�$�|b}�-�Q� �nҀ��`[�nҚ5Β*�`sz6��`{w��{�e�|�(� 2Ra�V�^~0�3�xkM"|���g�,jH�`K�#��g�,�%�=���#���_�&>�A��O��RS&�N�1]�h�6]�zٱ��v�{��D�f1��ef���ᚚ��܂f�F8�>�6���cp ^p*��0jedݖɋ�y=~*��:E��'!#R��}�YҾK}�x}9W��,��'�S�q,�������wwvpڪj��.��~~�M+���*�V��J�����X����1�_�Jg��#�P�S�D"NPWBϸ{��&I9'}N�Z�_��DN�����=۹75�E��X�E	�ã��o��M��/	w+���Oz8��X��'nw_�,?T4����@ҳ��%^`��@���-������V�����#eecf}���l�9��t��T����x��	�Ϥty��$77��F�[����Ҷ�2����[�⇗:�~o6N���$.]ힱ�t��&� ��v�񙛝��M�!9���AU��Wh(�~U:`�)w?���A����K(�"����F�+�	;�9ztfV�k� ���֚9"}�	=NRH�����V'�C'���)�����r!��{\�d�t]��g�|Ɖ�,���sU��j|������M�)N�\S�hXKW$���C�(ljk=��u�I7vxl��@���qi�<��%�������2U"
���03�A*��'�r)y��n�yV$g�0��gF�&��)*vmo�4�(N�����D4�i6F�=��|)�ȷ=�̄��]nأ��T��y4�o������o��g������56LY��z�3��'��\>p�"e���������yR����u�H�ǲ�P�1�����`�Y���o�|X��I.�,�5��O����/s��P\0�F(��D��^dqdw�,&D�z�`��C��� �h���q��~m��hO�BS��C���]g����,�45$���jғ&/E��s<}^M|	^�l�RZ�5ڭ�;Bw�$��	�޿�(�X���iNi��,�D��TN�!��8�#p�]�Ǫ�'�J�.t�&��]� 4:ofB<@���rȪ�����ϖ���6��A�Ӭ��0��Y�#q#���K�����x�s���w��~cc���@�+ �N[�vͦ���.u�9�ۘ{Hm��xH���(��v!�I<��!�"ծyRS��
2Ƚ���.@+�䂍@�d_d�P��t��
�M��-���Hq��Sخ�5f��@�Z<ՏWK�+G:k�ع���f�^�%va�J���$��9�Wᣱc��J��
a�p�)��/H�M�΢��|���X�X R�����՞ڗ6���Z`�G`�%���� 﫥D�OF�þ��k�}C�Pg휳}���w�<��� �RϾB~���J�pF�lM�z��w�^���9y7�u�D~g�J$S�EH&;�z�K}�6p�k&UD��Kb[c,t�/�~6�
��3�_�w���<">��0�[}���x���N�E��b/�����$ih��O��>���ϖ�����u�ik�%��߬nm�8�������p��NL�݈ryY��p�	�`-��{��HQ�C���y@Cx@n<���<�	ߗ|�@:/�D>�M+��C7����#����qH��A�3���z�>�����SV�����_��M�|�gr�Y8�iD�f<��p���@�D��ט�\e������썴]UX��|d�-D�p%b"X����k��D�������Rɪ���t�N}�����u�������V�x��u�n]5�|Yp�VF�8�܏'L��F������i�<>>�}-3���<��&��歧kN�Jwױ�2f�GSC�xJ��� �K�
���|M�lT>r���]�>�S�ߊO�J����w\A2c"�`��	�R3R}���f���`��UY���+��("N�W)��?_�*��
VK��֤
�5��[��\R;u��%=�q����ɹ2]Պ�q�F?Deܻ���מ.��ollB���w��G-^>Eʰ�8����H��t��{s$^������v�*���r��F��o�E�6��b;���$sڷ�sD��cߟ�bV�	��~_[�?��;'���ˑ�?��#ۥH��i}�[�`!���g�B	;r�TsF����`/'dff�~�IN�o�C9�ݱ�l��[-W0�WhO9ŕ)��_%�zqmm��t�y�n�R+x���#-8��u�N�V���D>qS8U�˒0�2�ɥѵ��4�/��[�l���NIc��$d�V������im!UUݕ�N��m��7��^H�]8����[U&�k�`�3���I�Pơ�0-���L2�nVœ�b��Α�O#�
(�nƶ*7m�#�O .���8݅�(��ڎ�VJ���U	����`kF�؃;oi bV�ɘ��{��+p�z_���"f��fi��h��\����yQq:�/uU���p���.Q�D���LW��J����,��_��U��E|$*��
���&��v�� l_��݄�FI	���v	��m�gW�8�� 5�q)�B�����bDMG�S���e`��t���ڍA�|3���������G�y�|��\.w��*ɮ~N��w���R}��}��A�W���\^������@��*�η �a8�������m(�\�;�d�nǑ�vaF�R�n�O�Z����h�M&d7C����ɓ��~aa�YY�i��p:.�3�S�D
q���6P��s�K��S���_�E+�Z����`e�/�/����!�yQ5��5�T\�A�撩4*��>%zIY�SUJO�����������%%%�R��t����T�M����"s��O>G�������."�t#]���HJ����K����(JJ	K/�t
H��.%)�t/���������Ν��<�ܹ���m��+ݜ�U*��ӤU�4��>/!d7���,s=������N=����D��s���%C��͏��P�CS��F��$!pw��N芧r���[+��������Y�v����D��[9����\�A�dmmWe����>����|��s��y�'��<�tg�y���N]��;ő'A��#��њ	�� �N�w�(%���(���TJ^S�����m��$ţ�ǔ��U#i���+�<{cs��r� żK� ��@�C����#V��E��i�F_�|���h�vF�}f�m/��L�~���%����<_��ff��g��9oծ������(� ���2���D`�CP	UR�)����kǴ���f�<� .�K���(3$nB#4 ��?9Ҕ �Y�<3^X_YK͓>�"A
��9x��M+ �%'�Ɉ��=k���ѐ��8G�6��q���m(Y�o
�a�� ����62:�M��xՆ�t{hӝ<"~�g�m��%��fXy
q�X�����lz��O�?��!�x)7h+�u*c:6�����SuU�'�#���;R�o���A�G� ��?t��H��6H9��ʳ�Wҭna����<�?��7J(.�կ�o���J :5~��?�Imy�˹q���.*!�Q$�������U�"la�;����a�u����͆RI����}5933��'��X����zza�W��-#M~���60d����2a�ZfO��5��W�?eWQ�dP��~�Ϩ���;9 I���QOn�H�G���w��z3�=���)������u2���'hUm���v;�-ak�����ηtg��aDћ��Br���k)��̵Y+Ƽ��,f���<u�$�'�,g� ��_t�اII#�]�xj���]��ah�t��A�%W�I�,�4 e�rU�Ҳr҅�V{O (Y8x��YrETP�3��2���q-�,|���W�`}ǧOҽܸ^
��D�ԩ�O��)&2�D|�p���?m�����⽹P��ĽO�=�8jc�?�
}��ocE:ٹ���G�ăc��ui;�ރ�#�k���Ԩ>�Շ��d��&�#�v�ф���|S{3�0��_�i����qEk���8�7=�$�ɕ� ��~�lb��q���$���ؘ�bE�B�Gd$2A��t�vw��*B�æWUQ;=��QaeWi�r��f��*�-P�C�v ��ƾ���6+y�=�b�hSr�-��T_q�_��squ����Q/d���A���K:ܮ Gr�N�7���X���]�{����6v�� ���v:���0��+S7�J��1�ʻ>Z��FrK�*z�|��8����_'ߗ5�w�"kt�aMlC��O��d��mxi>L��&B��Њ��?Z��C��=�� v�߻ᡷ-�~y�f�X�:k.^Iى���sI�G]�n���XG)�Zz��'���;NN�aE�'���}@x�D����"9(��(qp� D����4E�|K���bW������|�0.k.�Y~��^B�H��~�<�¨|�(H���ɣ��7�/��Ytէ*s̟�O��xƺ��+=�`33�A�י��|��6w��!�H��d}X%bz�]ߠ)9+aO�&]�
Ĉ��+�%^�����r��gB��&S
?l���S<~���[�^�?�@�d�|TPƜ�����4| ��*�!�s좭&D�U�����e	f�w
ǥ΍h.��4ުCުH�}%�妡R'���^z���.��	�_�I����D�z#���r�E7�W���{�)�\ �����3��R#9Vq���d`��B��|@�d�����AP߿�v?���IU�7Ӣ�h+��������3�Sv�F(w��y�f
��eh�kF�;��{��J�,_ҹ����%� ��&hfN)9������2E紧�*�ԃ��KJ����������HK���E9���O+�:i�wF	,M��$@P�f u�L��Z
;s����7�(�d�Y��y��a+�4�b����_��	P�a��~maى���Uf�=RaQK����U;GY�d����w��uH@ǉ�v�]��CY�T��-��4|�K�x��^1���۵�=�����WM�$��.M'(��I�U�����yyv�@��=�<M/�aPnq}�3�����Ig�}��ϟ�6���ĵ��{����;��J�����	��q,Z���+
3���h��i�ӺP�=��gl�*i��8x8Ƕ �����z&����H���Ŷ��b��TBDz��a�L����Ǚ
���k��x>�\�z.<������F[�,��Ǝ������b�YCw�V���c�������t��jE:�L�y�\U�?*r
x$Ɵz:%1c��:g?��>����=-�'���$tD��E��I�GO�$<��� �����p�2�"�Pܶ�X����p��/��m�_�����{�a2����Ј��?i��,�P���]�^`���ͫkj��-l%YDBL�k�YN����O���Ɏ����:dV�1��'C�#嘉M*�:�xc�Fۘ���04�2�"�M�iRۗ��'�]��|\ҟ�di�7�Ѹ��jt)�O���̢K�A��5�0��qҰ�Sp~k���/�<q���?���"bg���u�P�yWq��s!������o=&;�]`��J UB���^�O 6����Ğ���Eu����}����U��|������L+MM�i������ע�F��̃�[g���ʗ=�ҘWnKz@����s�RvK崽�'=�h�h7�~��������������qE`V���+�O!AS����A��q�".�����_r��<=�c0drSS��\T�F}'�-4�2�n�;�S�$��N7__Q�l�{����>���˦��*��]H����|�z��L�~Dr��X��̚8PB#�ý�s�A���0�|��+D� �L�3A�5���g��5�}aa�k� ����,/N���NY��J��+)V��6�!�;^��7�L�pXe��E�ǲtX��q�t|o�~�jH�V��"S���M�#R�C������v�V_����!�5���i"�$�瑀ω�1~�l��U�~�qC����B��x?%��٤	4�z����+׻/V�W.�S����g��{k�@J��ʠdg���ɐ��J;��pq�����|���m�т>@zk��e.ψrB˳ ��^V��	��� w�5yrR^(���	�����.���q,��������zl�̽�TE*47�|q��N|Ez��y����m)��e�k�X����R�>�91
�i[���ߜHqw0,�֧�|:����ߟ�<���B]���7�jb��S�I��-���R�8�k%O�;�6�=*�$y,IIh�4
� 8�*��K��r:3��(y��(�LF�F�����S����f�`�_�f�6�]���0�(��0(�??���a6�28��b}1��"��c�X�"�Ƣ9�x����V����n1]f��ͅ�Q1���7U��9�?�f]I��!^�E��^���D��e �����\�2^���	�	~@T��.�4��v�3I0Q�7�ka����0n�����9y��������q�ύr�B���+�Y仓�(F>+����zXbzdjj�	��L�*	����!X�G�/# w�K嗦H�����=@������:׿�V��l3T�e&��8J��:M����]}�I�Q�ۚ.Rbv�P�"_a��[z�lk	�i��|�$�%�R�{����[���Ӌ0�N�v�0�Q+�U#��l�*66v�ތ�V��fo��o'�]@���W9�K�R�����T��hN����>͡���U�w:��2�S���2�� =���Gl����R8�Ks�9����a��EQ��'�z��nP�7���]����+���e��~J����~��	+��@X*���b��̌j�#P��[��)rξY��L�˒py{�C����U�i)����5LZ�ꬋ��`^����M�=C�����ќS����2�/p�,�]�8��s>���i�k �2c�@R�oR��#s�����U�E�S�{�o�]�1c���
H�_��+�<��/�v�N#A��a�	��'���Rv��1�A��'�޺���]N�ԙ��U�t]|��� �NL�Tץ����������{�LE�j~��`F��7WL�	:Ó�X$����"[ת�k%)4�P���P9T���@��a4��OV��vi�Lu|;����t �?��պ��*c�d����~��܈���i= ����0A8�{�+ŻK���baqr0SA	�E�>O�?�:����%���o��_��) ��97U�D�T��!�������S.����W!�,,AA-���a��ʡ���-�s�����L�y�~	����5jS
��N�od��kMh�</�I��*Kj�Fk(�=�׫_2s~�|$�'��!�euZ����D@�=���;�� ?v���~Dnf���i9cy[ Y��239r�f�zv/��[�1��݁_�E��e��8
�
��K�7� �ER%q�"��}���Jo�nE�*�n����P���o$[�/�s�붖Fz��5�҂���r%kٔ���^U���h��v�$���{�/8��yl����KD��E&x�0c�بa���T64��W�P����8�L���A�ǫ����O!c6�O8 =���KO�Q�~��VwT��kw�;�m��	�N0c�z�Q>3E�p=@�u�#�f�}[ΰ������I�N���c@�)i%9��rty^�4��K@���V)��cwW��~��+ϻ��~�кO`��i����c�Ba5�O�"�����z绋��N���6B����jT�fNg8�W��[�k�A�W�߃C��8��"���c�l��F7{�X��I(�3�x����]Z���Y�Ã;L��2�@P
�5;�HM<�����x7�;y�9�c)��j�
�X?WQ86t.��\�~�~ �e Iw�P/zIpx�w�D������2������ȼZ3�#�+Dj�-���Q�D���ŭ�`_8�ց�%w_��'�>�`I���""Z��YP�e��췾'�=�ߣ�{�����07�yF�K�9������	E�Ng�Ӻ���^R���B�tk����7���Ӗ?5�7b<6�!���)Х��fu-gV���!�3�1�}�D9��PX�V'C&4@�O�V�D=
�r���a�S�a�X�V�$�ٜ��|�Za&�MJ��잼�~�?��M�\�~V��''i6�ٍ֭��Z�4���D����I�
�K�S0�S�S�%��Yxy�V�"+5�����&�I׻��쾂LjOAb})�y��q��>��C�Ahs_ޤR���}'�u��t�n�����@�7~$_��G��NF%��;�T}3_AW=�6��OW�L����z����R��}[����P��G}��'�޳W�y\s:��I�IO;7��4}'��᳾�7|�W؆�VR�e{1��Jw&�9W@#C���H��G� ����tjJ����c�֔��Ov�p���fn����T�=9����Z��R�`\/��y\�wH}�j?���U�N��%�@�y)���C6����w�T�\#+J�m�ɽ�K
4�������
�N��~�b'�ؿ3��M:� k=�Fퟔ2�[��J8�U`��k��o[]����Qv�z��vmhh��z��_�)Qh�: �����!IlL����߇�o��J��_1L8
��J��ޫL�̣�p�bX�s|a��Tq��AՎ���{��l,���ߧ��zi�W��''�PC���C����
ܭ��x!���o��s׳���?H�7{p;KCތ�RU�iKL�N�yw&!3h�d��%^MC� �?{#�֣L�y��t\����I�ҵ4�>�pQH���H���9�|�N� u�V#��Z�R~pdW�l���E'���������?�����F�=���hV-��I�X{�Ի�67��D�b�cV�\3&�+��~����>�ݙm-��q�]����a�I��x�576R����]~�/����CH��x2�~3 �	
��rv�e��|#U~���,��H��r|�>�@�#������++*,n�TG1��n�77�������
�ٖP\\�u��HK�,����Z'346�K��{P�T�C�N��;/.���3��Z׊���s�-�M�훭��r� �!�rd�0�ef��I\��]pӒ�b �n��#ŒGY���fN3S䍶�|��\�[{���c����
�~=O�������+N>��\,xdu��Z�Q�R��4���~��� �O9H6�+��?['i�3��Q"&Ǥ���z3H�cI	/�����3,�B�E��FH���tI�޶d���,A3S��.�T�/�e���x���UQ�ˉ�ç����ퟥ�9�~O�� �PYWgW������G���K�����o�������nN��}�1���Yh0�z�5�r^"x�9xy)�U:��S�uo!��S���C 姫'N�6N����Y��@uuV:�uR~(������X�����H&Y�_U�����o��"I�S��u�������4>�U�4ޔOv�N����9��1��[__oPs�tJ����m�t5(8�X$�g��9&>9'��K�!d^/��2��05��xX.���s9[������9��z����W�K��qo��c?��=���N8�������`�\ӁM�����rv���]���U�{ɪ���eѩ�0�A���E݌ȣ3�!�s��5o�W��-�P�^�1ˆW��� �wSk��h �h33���,my)�jSUE�cnBf�%aJϺX�����?>[�-6��y�j��q�$%5u���up��"��
d2��u*��1\�,��I��v�X���4�N���J��L��,L\:���t�O��m��-�_����,	;���R��F�u����kà(���iW��v���]����5܂Q�{;54�8\O��fw� \�U���듛��K���e�����_�������egd���p��*���,��I~_��y���ȸx�B�_`���}|0�0�l�F���<t� _�� ߢ��ak���!��n��u���S�g����LO��]W<ovM�H���W���x)gn�U]]m��Է��i�e�\�>�A��F��O��=�h�?Z-8|�}Ju����Vl.���V�C����.w1���5�>�;LF~�)i�_F�sٛ�3=}�r_:Y�Ԇ���who�>0���\Lpq��y��q��{�b	6�7� ]9���q���	*�~���+!�ĻS�j�Rm��ǘ�"��Y�D��r_�+P��X޸�?0_avј 4�0��������wB�>�݋���ܤ�̵����R�w%�픈�봪pH�;P"J����k~�Yq�M�f�h���"�i�JM�V�e$Hօ5Id��#@�]Igu�)@�n$:Z����㐬0ˁ��Q]�̂����U~��-َ�$J떿.VVO��7�1<j0��~�����-��Vr6�!�a�S��i/�~�5c�4f�/al,���"��⽼�	���j:�j�kT3���M�Mr*��<؊}f1��<$�U�~���jໍ��+s��8b��aW�E�V�6�6��u�R�=?2�x��M����C
�Emu�ѧ_���=%��3.ӯl�Y�l��B��4�ÄOH�Ŭ�u��[Qxs�*�XF�����I,<������,7ifO��T1�=N��F\�s�Ie��-,�����^�qz�	��䋪oP`��OSÑ�3�F�����&�dP��](KF�(���m�cg`ȹd8�v|�`:�7������q���^n�D���@rK!��>�8Y�ڥ8���7��q6r���Z��w9�������z~D"�h^ب�uʎ��ˍ�F}�_T���%3W5��>�q�Lv��
��7� �����ͺ�(��،���#QO)�!_��Fo��/ˮpN���z�Y�F��9d�_�����ir5�"�L*�}�!����bɨq�*WV�s���?0�]�N>2� s
�2�S�6�mM]��ߚ�:3s�'��	lD��S&v����Zf�P=���1�ۡ0�+u�ό�����r�;�˙t�ΣA�3#^Ϗ��OF����
����~
�N���I��D���`�?��	&p�H~	���}A���q�[�b��:y�.U�6���'
x���ׅ�~,��2+�h�@����XV�
�����y�% (}wqʁ����,IU�QH&��UDЯ��웤��Mp����(��X���o��(]]wث����⫊��(�R���G��>��a���i
��b�����o��2�Scs3��%>���<FBL�$�}�<6�ۛ)�����_+�$��h�JL�+mD5���w?Cw�lW.�F4mL}Q�?�~�8�>E9�G��6���(	9?cH|>��M�v�@�MAِSKuI��މ���c� A�T6��	���<weSv�/���Փ'�� �^��4��mZ��5#-�h�tP�-��o�ow`����ԄW�ⷢ߮z�W[��tX��$����vǫV��MLlz���n�F���V���R������Jl���h�d���[v�/u��o�i�]zV��K�@�̄	H�~�NX#cEA�ew~ff��kYk_`q��R�/�|�-<,��/P�EAi�Sp/�7uE�50�T9��M/�M5j!��R����bfH�Qc��pH��i(7e�!�� &S��˨hu��:B�qH[�0M�BYO��R��m�ST1�ԯ��HI�޸�ΐ+A'��O��	J\)�����`:���a�H�Ϋ���{�v���1'����s��a�8/nK,�{=/@��`�4f!����c��M�Y�"D�n�<vs�?8�?Ľ��� X�DM3�مE�39ʒA�_�vM���AU)_j�OX� nIE?�*'���������)ۈ�����y�ۍ��Fl��0-)z�cM��?�L����6q~A	K���W$'�A��T�լ;a6�N�s�[tV����xL���4��E�!��Sl<1��gݨ3��k���а��03z�q�D�̅��7��ք8}0�&:\�Y�eF,S:~������x&QrV7�.��zq�����ܬ(�eA>�"��#͐>�T#�i�HB5u#4�,�n�V�u�6�:�����/p���z�t!4#rG_����!�ɂ�~��z-�u��"� ~�a���r�/�Y�؀p�WElU:K��NھbR R�C,M���6`���<ڝ���j4D9�xjM���y��t�8�+!�l�m��5?�[�|�K��:�}����vzJ�����"fØ�F
��ϽI~ҳ)���y��b���3��0{�Y�WލT%�^�~%���m�����3{��H?�½� M�uN�!<Is�#7��JE! �(1�#奓@|�UݏN���k�'!�]�c�_��DQ<��<S[�|���d��Ӆz�j��J�C��$3Q��r�=���}�w_�EQ�}Ѡa��#��ݯ%//I0{�oH�����q
�v�:�?�t�"`����
௼��F�c9O���/���܃v0�h��x� ���j�]y34 �ϥ�α{	\V���SH�;!>#�,�N�|f�`Ԇ���8���^Պ��/�Y h�v��j+_T@��W)�
GuاoiL�?VCRA����G8x5�ix���M5��l���sNz���
~����>WN�-s.*f\vK���Ɠ�u���%%���b`+�o�- ��]HS�`d~��W����T���D��)el�h�gz��׽癛�?4�M:z{f����4�F���	}}�'�06��v�|��ڍ���z�N���F��^��*�a�mt&�S<�V 12��<�S�/�
}`��AF�8�35=@��b��P�H���
��O�dh"9A� ��hz���^�pE�#=P7I�٭�Yn9g��E	M�7�D���?��4��V-\�}�dH���_�=�
��l/A��|1�/����Î�i&P'�/�t�^��]:fw��^~�b:;���k����9�k�/�� �����^0tZ^����� "�#��i{�[��;���]J6J��O�(E�E���L�͏��Z5}���R�
Oo����l��p���i[y���I�c`�;��Q=$ƥN����ԛBPqbCK温�ow�H=@�zn�ޮ֨#�hs��@jx&IB&=�3�a�����}�X�*��ԭ�QRRo��C�t0���~�l%D���!9f�9�Z�3��a��w��2�nÈs?��)sw�:;-�Ћʉ�����y��v-��O����^����Qra��hhX��׳)���=r2��3V9�~��Ǟk�& �u!N���פ����I�MB��Lx�Wg����Y^��m�z|=G����n���(*��x����M 5��k��� _N�
���u���A��!PX��q� [���b�'٣��a��T9s��׍��9no:H��c'Γ�RFْ�l�����}���Ix��,������%a��ӯ�E;�hZ"���r��8ā`�I�tjv�����mI��
㲷>9�^V�]��SoY�.b.��Yj���l��>p0�>󇉀�)2���(��ӻ���^k�鱃Mj���d��� ���2���?�Ӷ�����Vr�{�C���;q�����g�9�;�_#�g�+KR�[�W�?�Y�����6"�$�Bd�Z�*�Ӭ~��@mo
��؄�֊��X���b���_����Y`B<�ă��FW�j����ꄸ1�)��̸kޱ��V��������h�}b�i,�5<O`�t{���ʐ당|�ԉ���)�i�\Y�Y�����]y����{���(�&�S��9���va��ڝ��x��	KKr���2�=�K�>�v���2T'��� 4G���T?�F��)�zq�M���VE��$�e�
F�_e�rUmi>��~o�pѩ2�$���A-�qߔ]Y)`a�/��L��'>��K�E��Ta�O��P��E!�2��'"y!@���L_��'���y(���'}����;9����؟�/;=���͵�e������8�B�`t�R
�wM�Z?[�U�v��W(�����F�W����@i��!��ay�[�����0=W��q�e\J���d�ȸ�a���WAo�q���G{g��R\c[�M^�>��@o�<�I<1^�`�ɺE:��n�����H�+��cE��֌w�ý��-Wq����V���{%3o�_�P+ao�����ݴQ1?r5$vss}~6�I������bo�z�G����q���_șJWJ�3����ย�GDj��BmS���+@�Q9l�KQ/"ԍ�.�ՙU8���b�5D� ^�"��w�1,���[{5��?VkC�n�Ţ�#��O���7������F�C���}U�҂�E1QM̽ny���C�l���O���%]�8�|��JW�ٹp��E�7������=���.^���my��=N��UQ�B�lTߖ��KcR�Xw�p1ԣ�A��.Ja����pzo#��i�&K��`d ���媟l�gGϭz`F��-�vwZ��b�_�'��k���5��'�fsw�2
�`-�w@��e�ט�$� ��͇��ݷ*J�Q4��l/܀�5ݛ�U�>�����z���t�������(��?�u�;"e	��qj���7(vS)�.��ʶ��:u�9�A%5S�P�bQo���ׁ������D`I�EupK�6���2���4�Jg[�l���*�Q�$������Z�ZiB*�r�91�iq7b�u0<�<�f2u�"uڱ�G;c0J�)hv�MGǙ�x(u�k�o�"mo�b{���n�!��L�gV�]��{A����(�~��p�K�}����S'�*B��4l���>G��.Ԇ�˷�k�E�t���m?m���E5?�S�e��S�[��_]	}y}�e_�jPgG�;����ț9�e]�N�3�'XI��@��Z��(U��Z37���SP6�DJ�8�\V��"=�$!D�CNL0.k��cO��툐?X�ϬCsJ�a���/#�E��݄l�l��vq��򉱘-zl;�LŪM�M�6׻��J�ڂ#��7��>�	V�p��-u��.�J O;p��k����ٛfx-�2o`s���n ^��ڹZ�ǯӀ�^eҕc��73����ڷ�J��r��2ɟ�|�J��?˙�Dg%��KWא���f��dG��3w:��*j,��r2i�E����]P�m�L���$�)KP&f���
@F�^��6CR���L�b�u��l�&|ѱ�V�� x{
"9D^��fG"d=�?�"w�a�&�G�%����Z��.]��mp���O^��=��Q �8��<�uN�؀}�2 l�+f#�m�:�ރ����J��3�2?IY��M�
���ne�/e�!˾ŝ�.84@aw� ������PVM����kO��^�/<d�N�5s�9N����e��O4�Dʹ���C�&�[y�D�@�[�(U3d�	)- ���wgb�A"����Л�o%�����>"������C5��]�N��b���ŇL����:(r�����%+j�,����SH-��_q�g����G�����m\�ƒ�H�tV:�5E���CP��X��c}��ƺQ�UyiA��an�ū#��+��R����u]* �{�: ��3cv2����bTء/�&�<�"�/eP#é	��+��UM2 �a�&�5�vb@�p�]�dB��MZ�)P��������2(��8���'E���T!['���f�ɪ'@I�X8`�{���@�t��A���[ǣ���o�9�	���f����X5�9�/f,/����]����f�J��Q|c ~��۰#< 6�pF�ӂۡ�I&r���ȇo�zxx�DL�Ɓ����*n�@�d/� (��5$��q�b��S����̤s�#�䝁�,��u�K��MB���-g����r�M���6�ۓM�p����7�S�hܦ��i�����g�1iN�fH���~�/�����LlaQ��L�.b n��B��i�UZ�0�i�_��~�V$�q��H]������EIxD\VXԣ����OJ���ǃu���dE"|�?wށ��[ZϢoR�����ֳs�i�7t7�	�-o48%�u����n�YH"�k�Gks7�6�~�)�� �jR���/�FP��ԓ�,��I���c��csĩߎ,}lo�yys�4s����4z��\tw��l>��6���+s{����$����A���!��ɱ���ܤ���9��zUX3�q�.�����_���n����o���2��S�Z-�L��,�%w�:+���O��S��BXi�;�����d2�P���t��X�R4��L�Q�/dL*�.[+�د׉k����n���g��&\ ��Z��-f,Mcv*��u9�l,ǩ"a �x���,��o���Lihii�|}�
�T�C��+U��RC�6d[���\GK� ����1+�f,wsiqY�[����	& �+l�
<�"-��9.b[m��[\��^m��lP�5v�$��;��'������U���M�����	-gK�W?U}�7��Z����BSO�Oa~�^���_�%�W
�[/���w
@���A�;l������>����6�y���S2�Ѽ5�Uv���ԓV���bh]7.Э3Ίy�?7�'��c��O��K:L�7;���,���� ( G��bo<����u~Ŀ�;����Ŋq{e�͙Ok~��avO�BK��yuKy���IɎu�s���A��Ϫ�G(��vC�f��#��a��L�^'�\p]	q�yk�����rצ��W=��s$W�jM�Rsӆ/��q�W����_�g���Gm��Ϗ�Zm�r3Œ�O�g������@���E�e� ����C�T5AT�"��@j�;�rx�qY� [�L��P��+00��u޷���-YdksKNj����,Utu_�>q|� 6��;Ώ�B��|yjFo+��*PR��o���82Nca�%���sF_�G:��#����rc,^��v��r���Q`�s�������]Di�����l��YV^A�#�����[�_-k1�@�{3��������(���;�ަ:}G���A���<ۅ*�N���~�D�+P�1@��o!�o�P�S�!��f��ld`R����ϛc�wv��]�5j����=�����E>r��b�&t֏�9i�[�>3_EQ�7_��46��ޫ��I\��F�Uߜe/����A��7���k�V�����S�Q��DkCC+���9�֫���`��������:����	����� ��5�����ǷA'�}�^�|{6��=�8D����d�,�ۣ��.::�����ͧf��c��v|糭�s�Yǝ��2�jtB�l���1Qr@s�]��'��焪�VA�ˤ��*N��A�r����hu�q�­s���EG6fj�꓏=c���n^CP�8��sٔS�����Y�;or?@k���@eOA��e}�'A��o���	���?����A��M���Q���-�2�m1]�n��Q���w�Z|u������͑�H;K��_��{�-8�J���Л��sް��wD)�!��'yo��Zi���
T�}�&����K2��.�܇����p���эq���������a�K�)un=5�Q}Ae�}p(�)ߘ�zĸ�Ɲ���UY�Y��T�5�C������8k��ě,�B	W_����=�����1^�~�U?�(�c{���7�:�L-~TGw��R��u���I����+#��d�T c6wa�e� A!vD���{@3����At�����ʟ����~�ũ�=ٓ!oU�ۛ�>�@�A��^��~���)u���O[N�8>@�6F��҃jbﵲ�������X����'�N>�X�����0�c���,���wCtV9��7��4j�v �_|Y}-tn����n*������v큸����V1a����G>v}�2bZ�G}�?˿����Ϯ�������0�N+�&Ű��҉*t}V���~�O3�Ker�����'@|=��V�矞��kL={O�Gh��%SdT׵�N>�yB	�0�`�v�����m�T��8�DԚm����S�_887���MU����F�o��!q���Zn�aN�e�@w8��[ҿ�����Y����R¨���vBo�%���yW D�!� �eQ*	�gi�Y��9���l��T��I�>O��EA��)��U����^��7�C����#[ǘ�Ҕ��{e��,`��rL�����t���Y�!"+�ɱ�� ���ڹMQL�B�k^�߁����5)T@`��n�8�'�7hZ�&�J��l����Lwd����r�H�{E⢽7���.�&s��K�;��폤A��=M�� r��H���Jhe^:���s}�A���J��e>M�I��E�P�^��gs���O���qv�`ߝ{��8�^5��z�@�D����nM��R�����z9��^�8�;�+��NǶ�)�2 ��5{Sk��9Tv��sӶ�=��[�B������nW�$��;�x��=�#8�Ы}����@�|�v7AVs̮W���C)�}�ؠ�����#���n����4r��$$�இ���?�k�R���A0/4Ͳ4�6E:� 9�p�fS����_z[母�&�;���R>>�ݱ�'�'j���6�E2���,o���H�Ɵ�O~;F\�_8��3|�8���^�`����ǽ����P�K#6'�r�7����a��а����o(���Rvo�w�02���Ĕ�2}7m�2����i�1b�qT�N�EO��{�gS9_���N�BdM~D�c�E��9��O�F���@|8X��>`j��k��jP�����+���a4n i& �4&�rs�z޳��̱\մ��>�ϱw�������wCYC%�����B��5�-�k�n���0T�ԥ��v ��}���I�߽���NR�M�k
�g�����:���t�X� E���^7'�r�L�f���8�{��wH�Y�q�P��mw߸�C��z[�ȿ�x���/%�Ma�CP���m`T���ז��1�O�A��/!������ 2���q����ivM�t~-%���#���i+�T���\ӿ{�a��kx��lnݐ�c�Q��n��q��ފ�_��b�,�L@B�F<8("�x��P��|,��}���ا���������`�M�IY��,��DN�X��4��E��.����*6sA�x�n�w�B��^��t���	�鬡ʲr�l��C^��*����ܜs;���l|@>���W7b�.�,l.����ZB5�p�z3x�ov���V�jZ��\�Z�<���ޖ�`�O�3�f��A���ֆ�f/�9��j��4��hNLv�$},���-����=��ٜ��k�Ǣ���L�tu�b��ih��ʷ��_���.Ao�%�*[�"Pe�+H��rߺ����U}�!�PO����Z�sV=���q���z��T*�L�Hk�%��hV����~g�.�����Y��L}uT����"�H
()R�A7̠��tw�tJw(J=)�� � �5��м3������`��9w�}�>����}�T2j͡Wf�\X����v2����1v:˥��y��F��\��䢒��#Th�)���a��F���:�������RX֪�$I�y����@���jB������YU�0q&��'%n,�&O�[�qm��YE}�:JUdX��*�|[z��k.�uk�0\�����"�x[���5�0tR#��CW�j�ʭ菊�	��t�'!pMdɭS3'}e�L����a�_~�v���O��ߠI�Y_.��z�i��������f�%���V���pw���:���Ҭ��u,Z�F�Ӹ�|��Y��!���60�L=Z{r(��ߒ�/��67��n=�x�V��4��e�+L��^���7�ݭ���A�o�F$�a�e�|�b�����28����m��>�榬�Qgǿ�Ԉ��Y Z�	�/��H�dE���dG��Չf>�Gc}�\	I�k[�?>�0�c^�R�?�0�%��
Mŝ��F���
;���Z�ɚIW	����]���S[UEw���[�:V{=�A|���f��:H���Ϸeav�XM'����|�3;$E��8j5�t���Q$����l���;-,Oz���(��ߏ+�7yR�_��r��(��=l�ϧ�:c�@ZA9���������b������骛���ֹJ���-�iV�e��k��gk�+�%�oht@��h�S������<�u:�n�q�[�u��߮7o�J���&��W�!�Xٙ��e/��
i�l�Lz��F�W7�y�������
�ឥY���	�_�[�*����5R\�p�f,I�b4�S�C��o��29�b�3�*죪�Ϩ��5n��T��P K]鋫�G/�S�]fb��䡿��gs`��ÏF�5Ė�<F�,�E��mN��� ˽� ��:������v`�]�_��� nR����ǿ ;6���?ΤčVٖ����e{�x\05�1gL�x*��Z�w4��c�m#�96D|hG�:fѲ�k8���mp��#j	D����ԛI�ߡ��EQ�ؘ�i�ո��=��Y���9�moI:�6dI*�ȁ�"O������(���'���Uq��7�/��#s�/�Ф�D�`[!g�肘�*�Ǽ�Y&n�,7�y7���Y��uhh�Ͻ��.������U+��=gF]c%5��|����䣦�ԁ�����x$K�[�6���cZ�Wώ�ל�<-)��|�٪a  +8h����`WD��ݿA��C��[��_�&ؒ�cx@�!���C��5b�/�@kX��Q�*��J}�ﵓ]��f�{���noq�U��;24����U�d��H�E<}���R]�]ޡ3��r]�%�4��^v�����X�Y������9���pr!����rB㫈C`@7�828Z%����y�1���]�2��ܙ��ӧ8��h�����	փOl�O��a��0�������I�g{�p���}	��V1���Cmƶ0�`�u��+�ž���]@MP���;�XO�\~���'�X�n�R����l����' i��^^�#�^�a�ZX"���	f# N��}��*!�X]}|t�"�z�*��f�N��1
]8�����FZ��/� ֨��`@t��A��������b|��HxL	n�S�Vd��e�%%%��t)B���en���/�F��=�4��'�f��A�#|Gw�i��(L|�~r֩}���N�5������槑�9�G�7�F���)>g��O��u[@I�k�7-���x��i�q��x����=�D]4mZE�����C�.�=���4L+�a���9
�6�P���W+�k���BEmDM���X�ؕpx�O��J{S+|LÎ��n���t)e����Yx��s�Rٲ��-���u���G�<T��Gއ�/��[�o�լҍ��1�u�o�2j�d��;�]?��t��k�H+�J'�z���B�0k��u�9��{Ew+3�b��3�m��I^O����@/;�ܶgl�!>�H�磔K��I�A^�(7��jQ�!;�&0���i�a�Z
m�nǅ�Zl��o`�Dg�f������p�z�U�"�O�k��%��Yg&[	b��٪a�����}T���ly'=��2�G�.��z�)�ߑ�1:+`|��tf��B؏m���ڣ#l'��&���l���A�,f"f���#�Uq�[�� \n��4�S�ssM>p��~BG�Py���Y�W~���\D���$����aQ�>�:L��(u.~.�N@������Tzr��<㋕�U{ʕ`ԧ�|?0��t~/��.Ռ:� 	��y�k��Z,��Z��w��D�0N��s)�=iB[.�S���J��1�V�sS�j��׊I��ϛ�!�[6��вz@�����&���7������� n[|���F�����6?��cG<_���Z'���6�(�^ǑD<�j�X�-|3
8����G�^\l"���w����_]���5]�Ȣ�!�c��|�$Jq�>%i��5��%7Eǝ15J��:i��$V= B�~���Hi��� l8��Yny&	w�e�΍'c�!�=�^&?B�"�mw�33�����i��s��g���%�2<�Wj�Z`u~���'�+D��-�q�4?��X��)�I���E-��i|�S%��+�r��`qs�P�vk} �J:�n��k�����[[�/��w�)�����9p�M�n��L�����2��WSl=	.~����&�(���>K[#�SO���]�q�<���L1	^rzg�"�țV|�Ӱ��#��'e�ʑ�?�K��u�a�ͤLҦ�8�7�����J���X�t��d0ʢT?�q�_$Ӊ��Kx�bRw��� ���&�N���G��tMW�<�5��U�;P��)F����b�*>&���il�cV2s���L;0��n�d%Qm�r������@�M��η,�4q��B�_~g�^\�	f��x�V���*�p�$���ʎ��Aq������/a�:�x׈gmEƔP���5�| Շs�̈Z$���zM	?�}y짧e�n���n�� ���HB��׹c^�]�*I�h5�.g[�Bwه��gu.��ivT����d<�0-�/�VuU ��C�?^����=?�'����'�[�����M�ͫ+������̒��{�nN�*A&��'������_�<s�l�}�K�M@A��o ���~�J��e�qB����^��=��y��M��ViB֝k�A���4��_���GS7�e円��<�>�>��{� !~1�H�`�_�(P�а9Υ�ٙ�9��t�J����n����B��è�o�TU��cu��Рgs���7]�QP�Q�訿�-���}g�����|�pSw�[W'�k-.�����I�瞦�.��G +�p�A�. �����}�oޛ �K�R�&���y<�����0kk��[/�D�*	-B@��0���>5�du���$�S~��/�*o��/5g�[�G��BhЭ�h�0�YJ?�tȲ����a�� ��U1qz0���D�$w�����<����.�]2Fy���_ZT�t�t�Au�Bg��oMS�q�������y��7���Zx��z�@��������νd�(�̼�pԢ�I�N�@��R���ɹّ���2�z�1w�2F�1z� �����	(M(���t�h=$�J�N�n�nad~�O����%h�����f7�B�ciQ�y}�adEr0��b��1]�؋�����D|�{[��$���*U6�rs��\#M�BA2C�c�o�\V:v�m�ў&IJJ�� zܔv`Z��j���;�y~��:H�S�ȍ8)=�n�5�q8&4�s��Y�?|w�+K�����ϝ*�V
���:�I�ѡa��F��'��%Z�"��,YY $Ȼ�'r�6�(�G��B���)�f�zv_Jό���w;�������F��%�ЗB�.-2���kNCQ��q
�_	'U���UA77O����8>TyOm�*���S֗��jA�P��-0��Z�F����QNH����\�ék��~��D��6��S��~ܳ�H�����0�p�,@��]$!y�O���R^��%�X3Et�X�l��XԞ��^9͞P*.��o����6o���<iR�4����o}�密2���1�B �-o��|үыjHb��A�T����c��]/�Y!��op�4��rE	k�I���\Ć�2S`���D5����$/��'����/�B�{M>����B����g�W$z�l
BD$8�1�:�Z�=��o���l�u�P��f��!9:�q���?_u���B-�mΛ��L|I�ܠo>��( �����4*���&TZ>�K��4�My�Īc��g�ʻ�xJ$~a������C������aBD�`כs��N���B��L2�y{VIT�,����t������eG�	JV#9
*�a�hG=�*��!�j�qs������-�!ۓ�wH�|wO�
5,Zd�6
&0~����ʅ�S
\��9_�?�&X������<w��uKM�6ۃ�=g��7j��ҝ�M$ 4V�4�F�D���[���Q�6t��'���\W�����;j����ѐ��wc�پP�׾O�8��MB#��J��f�j�j5dy�G��9˝f�س[��=��rݝ��HY�E�rt~��5�J���*1?G4_:*����������p���<��,�ou��Y��*\ �4!"vp�W��&��8#�V��(fm��l=%�~�PK��v����K��D�0{����ie�ת�<���eb����f �H��]��7e���g����GB��h����g�-Iƍ��[T�]�x�@[�R[�W����Sǻ�MoZ�&�7.�����N\�b�êUw�c=�rT��H��o��pKM�$!��ɲ�@��L/�ebv������-z�e� դ�!�J=�{qAq	X}4�Z��O���NDp�?���o�:bj~Ȑw�0��9[A<���fY��dY4�Ӕ#�zb��P�ypV�y�#a�̏��J��x��;����?k��I��R?/���ލ�POc��2T��=�&���9�)j<�1;�tj ��N�?���/�X�t?LR�y��7C_c������z�ʹp��L�ʌ�Ț������~�����C3ϺCe\ˁ`sn%u�xL�n�����Dx�fQ�};p��k��K�j������)1u��E[�����;��)��Zx����^�<�ѐ��E�kv+=S�q���d1�=a�ng�28�0�����	���8��>5���a�&�qL�.��7ޟpӵP(��3ӥ?+T<W�B��6)x9u��H�CK���°�u�6ܽ	��z�����+5�����>*[�ʾ��
���%��g1���y��s��%U�����<��Q�V��(�{~6wx��dόώ2��^[&s����C�Ky,��|p�����7?,Rˬ�g<m�gF��������n)�9h%�� q��_nU�66y���� �U�޻��е��93|��]>�A6O1͎�n�9e�Q��ez<އ��OE��3�kAXXT�o�2��9�~�OǸJ��W�{oy�N�KSML�!؉b=}��S���KE���џ��@�gȚR=n@�x�����]��{�{Κ��A,�>�&s��� ��O�7;�}��\����<��,��ȉ����D�j��9�x㣧��i����h\�����u"a��� �(��V��R�������1�.n�� @c�}?c���H����@ �������(�l>B��bPq��lg�툱+�8�����)K�R=�'9��K߅���wZ�B���T����J�>�xy71"��w11̂�7>�~$^_��j�BG4w��3��*RE�|ӈ�
���>�χH��b���^�Ւh��`��M�PQh���@�]ԗ��G�p5�p	�$y�D����sx75�P�(9!s�:P�|N%j;�@��|��,Dx�Ӏl��u~L�?�p�T�3Y���/V
��q����뾝X�Ϋ��exϸY�� �R'aQ�;;�Bl�&���g���6��,�۞�TSB���G�:wE=��i�����,�`ؐ�T,�#ۯ{�8���d����\>���ج�Up�b��>�ي��ؾ�)�38�w~V�GM,Q�=���S�.��um�Xvi_~�;`y�R����x@>�z---�!L����9��:@&W���r������O�i����t��Yg���E�AC���RNyN�.���Z�lY�][��aZE�!V��2$R2fJ���2�%��yC�
J����w]���sEP(	
Ձ�ɻb�J�a�q��zP���-Ň|��� ��;��Ѻ*�"�^���Fk���f� 
d��	�z9s�F(�\\\�"����PBv1(�=i���<�[['���h��X?!�`�a�<�nXn�?�+��gI�ob�ɲ�	Lg�Y6�����k��s�N7���6sc������+�v^n��!��"�������K�����F���	�����H.,$us�'���$��y-�$9��z/���t�u��e�K��,2�GZb�jn�_5���sRF�?X�ϟ����fR�;�*�L8�_Г>�w�\����ͩRx�pM��)��0h���]�<Y�B�N)0e>�� �sq�Cn&���b��9j�k�9���&,ӓŶu���#�?�Z�?)��P�+K�w�j�v����|�Y�Uk���:	��A4�]���2r(g� ���~�1;˩����)z�p�N̅�U4�=|��#�Ȍ�V��9)K.Ki�o�j��bS�����)��-���و��ʉk��lnŮ�[p.���)�T��ц:@���O��]@c��Y����������V�]*��-��8�)�Tio��K\�0���!�������}E��w��=�j"�W]�������?�<�y�(G�S})���9��6�&>Z\������&��J{=be\s����:Gs�X'{�F�^Nϥ���\�V�~=g<��w��}�����]��	F�Z�(Jם��"�c8)��w�Gq�.��۷fmEOWH\��5��<Dx��K���id�i�`v0ȐH~�����?��^k�fu?;�������5��;z�9��b��\����Ms�w��;N����Q���F���Z7�Nm1.�88m��E��ǭ�p� ��z\?N��csmqX��<���pԬG7�.
?��3�3�!/gý��F�)6<�B,����:�:�%���6��4;o~�q{۵|�����='�]e.�����[/B���F�����+�7�W����D��8z~��P�<"F�{r�E�L�^���?��,�"B[V��M���k{�Q|_v>�4�=Y
ן��K_2���G���⠹�����}�$�<�9NgrҜ>�|*[�8ⱗ���\����h��Y󉵰�BK{,�z
���\�����{X7�z�A��9G�-wU�)zF�֪����[���VG��n}�efu�Ё�;(��B��!r׹-���հ�\��s�+:!�,�*V��Z�N%����qxo
�hJ4�����z���L.���8]juGM��ŮL��Le�y;� O'J����~\�-�y҄�*kZ��XsXY�g���=��_dJ��i�E
�������<��6�r����r��T7xQPNFf�Ƕx��k�y|�~\>�{�%�}��9r���}t���V�413�;�Vvo/;��Ȉ|�	vV���Dma�	?�,�-pk��3)**�\�Wr�I�#U܋�{�Y0�GQ�K[[[?�>I�������j�Uk�m|�`��#ח�f ��q��]�ⶦ	��Z����t��_�IJ���#z����J�۶Y���� ���%w	0X[q��ȄSF��ԳW�"��x�'�
v���������{�w�4�x�t���Z+猴ܳF�}cw{r<�V�*3��`�h8����W��ӵh���sW�k�-��M=���Zv�+$�NR����j�rA�	Loc��
�Ə����(�;����D}���3k�Y�
kMp1�NY=llB^Sy�Ū4�en�E)���A��Ҩ�}�	q�kY���E��N]Lk�X�l$s�.<8::��(����=���K�C�������q��tT9M�"�*��1aĈ���G1/.|�cɩ&��kcm�[�X5�F���7p��+��\��t����7:oȟS�?T]n���'
(y����5�d4����ܖ��C�y���g�%��Gh� 6�2,k��۳����)��nذSF��K�x��,��H��\�� �.�l{�	��p���H�R�~n�����rlIRNG1h�7�sb�+��uH{���I��v� �de�`T���j�6n�����Ȥ��7_�܆4oA;Nw9���Wz܄��g�ٚK�Ӽ���y�Bu���e�$G�^4.�"��."b�%B��:������S�ݯIVs̽�iim�Ĝ��bBk�"[��O�1��o1�I�{�����aHwq��s|��-sG@�3�e����cL�����Q��05��u���N��.#P���3:{�����L<*����2zhХ߼N��!�F���\����x]����ɇ�|�A��Lm����cqB�V��bd�є�<$����$m�I���d?'����&���"j���`��1����OQ�K�`��\���%��M����s4���Ǥ���4Vc�ǵ--���r�+�Q�z��d���wA`�Ne@(�7ȑѡ���(۟%u������KZ'����Z~f��R��较B�x�s}�c�s�k�"wj7�J_Ǧ���.��/�kI��STId&|���9��u�J���f��\B�T���v�J�DAþ�yƤ��j� N&�ŝ�^j��NO��p�(w�{���tَ3^RCx!�������U��t� ���q�'�X �2p$���~��ӆhU�R��Ɛ*�O�efZ�t�W����i�4꨼=i��b��@k8�E"?���=<�*o$�N4��n{s��Q�mM���K����v�ræh����d3U��.�J�Y��A �aB�/�;�9t*�c��էMLW_���Z�@��n�95!*r��D]mm�|L:8�h��V�o�������-��~h���$�V�}���͌ڄ������ח!A%Y�1qH��"��rЫ��gl��S��Rp'���8FhI_ɍ����#���H����Y�׋���8�L0&��q��G�B���u�L�D���u(�������5~���7V*N{<���*I����8)J��4�r?ܶ�bL�IEY�W��woV�����]\Ȋf:E{8B���,8&D���݃�7�,��D����o�~����)u[.�)�c�M��4�K��"zB����:H�4YЋ4ϲ`N�����t����ͯݖ~*�z�<b��5�J��ɖ6��-��/RA��,��g��tw��d���o���S�L{e��������]��ZIp�<�&u�r[���Z��y�ڿϘ�
&�~��Q� ���.�۝2B�{�\��� ֖G��%u~��@�lrÞ���XI���×&qbP-��A��������V�(��[ac��p�+�"�ֱ$X�.�+>���)60�r�c����j�V�l{�Ԋ�$ ��<>�q�s#��:� �ͬ=�!����m�8���c�߬��_���?�t�#��j���~a����^��гB��;�i��v��?z�x#�ECM³syL���m%�C^��u��B�?���O>���Ů	W��0��n�E�wH��_f�t��
���.��>C�6���M^9dW�b�L�Ѭl��F���<N�܃�(�El�'bca?��a#	�"^5M�8ڥ�����8_�nv��E���!���7���l3����kK]�q���y Jje!��f�/���=����u�Y��"���#�F(ϲN��g�``�FX�"�A���|��孖��J�v���0�I��B��i���'}x�gX��E���h4ѡ�j�E���4o�O�rz��{�������@���r�3Q�)5Q m�ʊE�W�{3�V��[0Gq��0ԕ�a�R��̓
N����q';R�U�~g쫃C6f�GHG;��(�����Q�~W�.)�p����?_h�O~���E���`�3��ˎ���Q~1x��=~����$HLg#��zܞ��]�F�q������h����tꤨ"���^!2�7M�%1$�Y�Fʔ2š�����z��s��uB�}���6��qf�o�����:IDt��D�x��l��2_"���FV��*�����7�o��z�d�d_���j.�d���I$���"���?��J&�]����ڲ���uXGJ��j}��:&�ydV��6�QuM���Gx��BC�=l��(���-��hS��2���9�yD�̆�6I�͚�4���| ��P�ըOW�D�5��ߕ��OT	���Q�]�GW�悒�N�0�^hŽ���9����^�'!�������B�~oV[n���?g��*><��q~gE��ҥ�1{�WW�T�<�@+��ot�
�|��I2G[��Z���d�Li	G���c�:
'
3';���Z�$�>x�V�;�����| ����\h��lڞ�6D�9����R�����=ȎS77��e�jq2�Of��p��ޯ���;�d���o4}���K���G"�M�3.�{�a����=z�����F��}����8I������j�h�Ar䍻�����KS�Ompk���W��Ï��D6[�%ade���Q_���lZu1��E���]�l�����w��
��a1��؜C{k;�v���J}��Y��_ǡX�ѯw�$�����d�ū��B��g{��J|ۀ0���o�}QϜi3���Jo��a��!N��r�JD�DKR�|����V���Bq�D�Yֳ�jɚ'>����	iY��K�R0X����d��~|R�+��ڿO�%|��s���}ٚ=��y� �?��G�c�i������X�(M�p�e�f.{ؗ��(�ٰt��><_���]1,!0(����� �X��ٓA����?�Ur�=O������Wz5�nz�z.�@��v�5�]!�a	˗4��N�2��)JN��RO]TdO~�>\�A|�so�����4��Mq��,^��]8�>΢�f�����ǂ�$��s�E|�zm'�0�S�]4��g��7��@������l�K�ċt�'�v��ݶrd#��j.J��a�bv7���+��sr8��	u�����ڸ���1���y~@U����\6'ɏ�� ����Cw�s���0��5S�K�(yv�o�ML�}j)����e��+UAn�맫�ǜM�+[F��!;k������6*؟�`�p��B�L��*W��+�&��p�ϯ_�C�*����Tq��ClMt��-e�kϤS��1\T[fwgtu�c�GH�"�J�(:�C7���T��W${$�y���h���A(k�h�rB﮶f�A���矍Q�¨O%�a�1sa���`���c����?�um>��9\��;E��J��*�Ԅ�2� a٦��)R�'
k$v����e/��u��62r�"��P�:�Vs�	�FG$2QQ�Y�i�yr�BU$E:!��Q|f���:]|����s��f�����q���}�u|����,C������}zU�s	�\��9��m/J|*�����j��(6|���e�_�����Q��U�ϸ1O������_��Z�t�M����7��X"+�CR����s7�c,|�t�*�"�^���ǽ��X�K��l{�|8W���i�`��?6�rP6�u�c�6C-�?���7�.��υ!C��vm��	�B9sp�Z�b�q�'��� �����!�+�ytH;|l��*���һ�4)�N�w�ӱR'	����[���(ɛ�����z�K�O��?�@�`�t����'����>U�Sy]8{�ˍ�X@Y�]��ׇTmΰڊ�/�ܝE�y<s�Fv��c�=���)��- ^��9�b�e�� Y;��3�u�?u����|�(1s��<]t��Yg��_�i�O�]KV�,��"��7*d�5�?�o�Z�"C�{Mf�+�US��٧dh:��(ج����XA>����,�7���م�?TeN�I�G;_*!@\QKi,؇-7�l���w��ͦ��q�[H��u�P)��Y� �d�d�� �0�L�=�d�Ȟ��m�8�����r���~b���!!2���=������_�+!�g���oy�92~})����M��<�^F/�b.37������	������9�a����#Ł� m��Ϊ�(�E�8D\�S�U.��*����mۘ��т��N�$u�����ع3�y�P6@���)��om��ϫS�d���Hѕ�8�W��T����u��q�iw�U�QD�u-g������!�໷'&�����$t�g�~�r�l`S��w�f$�p
J3�F�g�녀�H�c�G������v^{���-n����rm`�������t��)s�쬎��xAL&��a�N���0>��̯������p���nVgK�t��%#D���Ƿ^_v����h�����/�J-�s���#�|r��X�{w����.��1��͟�h�W��z���e�d��M૸��]�uc�
�ɔ��Vp��u���֒���ЧJ�eɳ�h�������'���u;�0����Q�V���ΰ��	J�a[w������u��<ʱ�Sq�ʩ��(4"+����wg�DRl����U�`�;e���k�{���x�l�{�I���I'듨q;3_��7����鱒��4�(���j������!{=������%s`��KTug��-�{Rњ(�����p�=�����K�pX���j�qWA������&��Џ��Ct֫�~������h�<�s��9� �H�H.cnV��>.!� � {	7ec,Ó���al@�3'��R܉�;��������E,�b!"��X�ɛ���\-�o�j��Z������=<J���I] y����!YcG����9Ӳ_�ON�a [>V�X�L���+!��=�	�(U�:�p0�;CW�Ҫ��mz����V�n�(�7&����v���{Q����u�D�1�Cs���w��(O�C�c�^A�չ����?��;+7w�\�7oBE���\)�D��2%�s��n�5�A1�l��:
YZxA���c�Ղ<��7���ڊ�w��C�T�5����v^'�d�+l�]%O�sS��ս�P�ި90J����طB�N,�h�vɳ��K��L0�<�~u�>��y_@ό�5��$�����%���+4]�Ⱦ�݃R!��F���Ӿ�\�wD������6�����]�/�����17d�E� u������s����Ƀ���Ҽ�읍rJU�H"����1r+�ą(�8d���m������c$��͖+����D�¾��R�T�2����[�u݆+�LN�H�L��Jr�W�y�+���>&�gVZ}%?�>�z�\Dn`�N�2����!��A#��3���G����\�q�/��v�J�J�p������zȶ���u'�i�������Q��a�������j�z�u��}'�J]��l����[
YZr{m�+�]�h4r3U6ڱw2y�vny���	�Ő��X7֌p�<�����o�!{�r�tn��9X�`5���Qkv&)Y�����XA��: y?�A�o�,�,�3y7��1tE(�U\OM�E�[A�^
n,�����M�K�(>�P�Fz���Z�鋮y͏��5Lǘ�Z�8���T)7Y����O}%����F�60�_�3���V9��skS����g�m�D37f�-qmB��"ĆZ��_���.��"z����%랥Yi�.��^Ail�a����F}��իv���\;1v�e��L��o�!����Q��v��y��d筕�7�z?~y��&<|�{������Mw0��	$����M���Ȯj`_믁��FA�k�����3t�OA���e�(�w�;]y�Ӕ��c��{`692}���D]� J��,	 �DX˹3�f���9��N{f`�䌾>��-�������F�Ǒۻͧ)�{-±Q �����Z;+��rW����o�g�R��Nv���s� ��YK��A��w�*׫�����D?6��S�H��{��{�%d{+;��z9��m�t��U�jd��������-��K2'�����ٚ�p-]�nİ�����.C��㸯�6<�_=3�?O��Z���ע��ڕ*Œ�
=ht��r�-�m�w�p}�p��z-�p�CWeJ�j�B�����d`����ܓ��:qC]ݟ3[�����X�e4�o�oG^_ӓ�� ��s1-xݰӐ:pxprJ�� R�0�F��*%�q{�{�S�����uh}g�Zn��{g�O>6�hiߓ/��~�0\!�96c}i�������*�	�LW���t�?B�z��;q�Ĉ��~݀��\|4%�5���Y:�vԧ��s�Β�E���^��U�[ݐs,���>���v��@aY03@e��4U/�y��j��jb ��r&_�o�~v���|���*`�᪖�}��BV5�ǤK@�+��k�����58' � �9����d��pF8)�_�_'_�Zε��-�A����s�Ng��^b�O��Ԙ��^o__���lM�4\ː���M�D{��5��z��L�Z��^�����n]�O�{�}��`o�L$����5�`�W����E�H�G�?��z	e����|�(�h��	����(>cuG�HoQd?�A�����n�+���\C������������v��n���Y`�۟f���W�ep�'�RÒ�
j��>j�{b���f 
�U���N�Sb���Q<�T���@�k���F�QƧo�/�;��z�Q[P��j�&�>6ӽ	�A+��e]@O.N�h��` 
y����������p�� �ba6����%�ݔ��4��/E�ޚ�
�z��"���5���WjL2�˛ϊ��d5��\Dx��˂��a��1G�B{������T�H��j<��0�8D���4C��@�Ã�/���9�쥯��1����z�����q�%#�m���̜g\��:İʦVQӛ���w�*�%�	�Ś��ry yS�J��xD[J�^���Z����Kv��n���"�[=*�;��Sc�W����k9���~K��^�0k�O��ռ���1'��1�ҟ��Ő�J׬�l��k�ix�=:8�ŏ�_y|��&E�L,����(i]Ŝ�kߖ�䥩�ܶ�6s������;�� ���x�0��/������y��B�l����:�ɆQ=�Ō�f0w���,wm�"�r�)r�ss�KU%����!U�?�����_���zQR�L0�v�s{w�uڻ�%����������]D�jY��5m���Q�/�^�D�����(��>��S��ˠC��:V��]��e0m�,Y24R�#�㔉b��F�����h�G�yO
RD)����1�^��ॕ���k��.ׯm}���H����_�/"bQxm�JMIᗒ�nk�c���446q'L��1Ȓ��FΫ4�`��j1����+�S���Oa�L�M���P�Q���/���0�������R-U.!j���/E2����{�x�5%�`f3S܄��u��L���͛�<t��ggg�|���4V���]�t5T��!�k�A�νϝMv��u_)v��^���~>goP!܁JYu�(�)����[@=7�~�;f�s>��bv$��}��Ȕz�?�^�G|���#lT����X������1!b�U)D��ƛ݆�hE�0$�>�X�4Q\y�x�\���Y������ޜ0sC^(<(��˲~�n�FS��S��G+O�4;�{E�E���Y׃���"R�Y�ec����`��_�K�fu��Z�H�)R=�s�M������#����r��U�]3\sv�秳��z��إ
���-T�-���~��� 5L��[�o��/�����<�I�OGd���(�].xܺy?F��;��m�02�G��-�oaoA�Ӂ���w�ߍ�+#�n�����-"���]M��&|��!ZvhR�
[.^r'���N��Қ�����Qi� �^�������s��Wt}h9�Ӷ6�k�� <�#��3ٸh��������%�}5d LR�q���������r��o}*��W,\��:q�?�vK�$j�3v�9����"Q��_#�|a!��t��9��
�U{��_TT���,��~b�7���ˆ.;3����:h$�B�����tb>ӭv��vfS3��C2�P!�!���XqK��r:��7-Q[�/o9*�"w��ܝ3b'5R�����K�cm�5���9�_��:˄ֈӃu�3��u��~d&�rl|�`�b����Z��mKrwM�d��F,����mί�:�Z��-*�c������=O��ҟl��n5G&���k�O�i0ƕگo�R�����j]�fn��+�D�`��D��O�7��No�j�>�Mi���c��~���P�,{$�$G�Ǌ��lG�
��������Q�&78{�P�q��͝��{_���~���ǽ_���9^����K��k�r�R� 4F@�
�q�c6���e��j���`@�A��/�d Y�㈆�4x
�'_f�����+��ѷ��R���ܑԢr�Z-.���6ǻZ�w^j�+|�bjsg�I�� +"��٠1qgh~Y_$��w��=�lj>:#x�i�3����p�����
a=r����awF�!P�٢��Bi+��x�bd�z#`B�\t�X��U&?:m��djju�"�t�w��Uϭ� B������S�OvF���rNk+/oA,��o�7{�AU��v=F�)٘8>)��Wy�'"���W��eQ���6�堜&0��("����k�'�^=����m��^N�`�5��t.�ez�0}� �:�1�:��vM��q�`l?�z�3&���b
z27;�U�~�"t������wL7�	?c5��h�Ey�5���]�5�ps�q�[C�7�z-88�{@`��N��()��F,qᛰ_p�&�f��t����F?p�)۬�v^��%N�
.*���@=%���<��b[�C��w���(��[Q����ۃ{��8����5�nL}����ks��ppt[�U&�߇"BF�O:vUPg�	����m}
�=xx
��M߹���Y�0�{�]w�����'�@�xi%��^���3�>G��m[�\��6���������xT8cUd5"0)���OS�P��`OvΎ�����ي�56O��|x���9�Q��+bW��.�c�Z}����Ib���N۞��牄�y�U�RW�D���Ү�-�L��ɺ�67&	�
BwM��f�P�K#;�K#^T�.ff橄�׎yE���m붌���L�L�sH��;���Ҫ�G|�K��\���kB�M��j��/� �c%��͡���|�Z|�c�f�G�e)�<��p�������� ���[�%�r ��&��K|�tPI:�j9��}w�7���kH�{������ĕe���8AO��%}��x:�DRR�g��v��K�e��%4v-������(4>z\�#���r�bp���q���?�?2��cʭ;w�K�t���p>:F���ɪ)��4aq��G�D�/"JEg�F�5�`1O��u����2ɼh�\v���9_��
jw�,d\q�U�n��;� ˙)��CL��ΜivKл~����(�2x{,�<c�r�de�c����|��K?�M�f�S�l!����I�����х���_�U��N��~\)N0*e/#�}G���}���]�"Y�u��5�rR\�	l�u�ǡN�j?�5ߛę �`cs��U���xK���3�h���)/B&H��昂&A�NU�	��z�6��)��Y���X���JF��N�_*��Av%??���_1A�ߺkP�X�Y�]�*ZhR=����;�|S��EsƢ�8[���]�hp3�̯��f8S�Z'CW~��X`����fDF�����y��:?�#y�^�L�F�L�ɒ�~B���?�<����m�3Xkc�]6x�}v��' �:L�q�,�M7��^�*±�����)�mb�A��W
ȹ��0�(����Oޗ#��s�J������#Z�`z���A;�<6~�)F�*��ڜ�����$� �v���L/Ek�!e�Ҩ.{��ٷq_�B����	qa)|6�`ft�:iO�}�'%~>���� E����ű3�+���<����WY@��O�>��6.�Oz�7�H_��}��^��{�w[$����ڟ^�Vq�u��_�I�R�DF���kE��CQh|�����QL܃���(c>�B	s���+������ ^����܇Z��~�~4���S{`�E�(�#*t�Q��ʢ���^&�y���d#��El<
�i��xG�/�Z�0&b�_{�����U�1���h;�#&m{J-�Aޟ�,�M£�C��J.Z�1Ny
�8s��$5՞�@ϲ�]˅T������Ś�����(�V�ᜮOw������s`����|�n|~��7�`�8����cR���U����^j0_Z�TRZ��un����H�
���S��҆�k�)xa}H?OZ����f*��67 �ޙ.�B{y��x��r���:Ϗ>p`�!��:o�L��:����*QK�w�h�����[�_-q��U�!�HR�W� ��C�0޽�3���?�xN�4��.�����35�� 32�Ѝ��O�8�)�$NGV�\@�5����U������5�^�k����,��ٷ��~ʘ�5J[/��27&0��ǥ2��ON�+X��g=92B"¾s褂(�>^`�r��*Z���ǚ�|������$�ӨL�K%𶼾B���"�U�.�3�b4��tKw�Z�N�򭩈?������<�v�4���`���qm�Qz�\��z�����w�6kc����z;y���L�-���.��'KL�Ψ�8f��Y��Z�k��*6��������.����;��AmRW�3/58��O���q��$���V��&1q
$iM�W2�R0��V��1
���,>@��Z�s����g�/��E�·�*���=J(g?���#=b���)VJ����ˈ�z�nP��;��zqO�����U�������z����_(��1�٭�_�:O������?��t�3(�PB��.�?�@T�HD�&2c��R䂞R�*|~&�)��*h�\����߽�<�<"6T�����[}6M�E�`g����:`ܱg��9�ò�,�m7��ŔlP����u~7]$��L�<,����3!�BSZ���0r6�5�)�L7H�!:T��������gTA�P���CËY:�_
�Ҏ������x]�����,��)�/���WN~+~�+�$7�&�wvH$d)�̍�^�^��U�b]��&�p+����b��j]�v_S�,��=������"�K+����H�{<�l�ȳ��2�GS|ɫG�E��ڦ�k�nP���YlL����c%��޻TO�2����U �������J&�x�q���4;;c'���m�U?0�	�?A/m,���
'����
&æF�^��K���,���I��˅9|�#ٰm՗xȉ�=�J\�4�V�h���)�u�|�o��q�0��W��K���ޕ?Ыҷ�v�5�թj�u� c�b�6��^��_6��>�떨he�/Q��u��20:��.؟�[���o��qx�T���uP�#vǯt�Urs�B��X�n������<|��g��V���z���jp����/�� ��"� �͉_�Z�����H\���=U)#P����~Y��>��ű��n.m��i������c~aP�>T~�����"&D$C	hM�gS-	��%WG;��t�z����<K��*����y��������~4ӿ�W0���\B9��u�Wv�JDH���.n%�f)Bq�pw5�+��[�!��I�^�/�v$�o�ؒ��	�&ؤ�lT�C�8-��^�{`f�v��p�\��i4�d��z���\�d�����rt0�:/s�����!nY�G~���OJ��@ Y���{���L,>�b4+�������X�%b���>1�rD����%Te�ٽ������{
445模��/�C��L��R<��,*��)�%�u�%p�%�b�����:����A�I knOxnv+W�ݠ�<��;		r���v�ZdLV'i}n;�e���V����[$�F��Jˎ�l�q��e�LH`E����b���W,�x'L��[Ak�xy:����Z��n�⋾��Wz��f*�!�f)��t�c�����ܫ*9ε�]gˤf25ă�c��h/mK�{<�{��'��9�Z��:�9�:^{�솿0�$'MCIi���G��|&�8s���b>����l�޿�4�*#XJ��0���\uF#��=�[.�ӼW����ٜ�_y���c!0	��:��&��C�f����4�_:�����R�Q�!/0|&~��j�^ �K\z(��Ԓ���E)9E�?~3���*QK�P�E�.�3�/�2��`8��-�#9E�Kz~�g�� iIڮ�f��-��Wb
�uS�vj�
�XkO�X'ݻ����?�#��	 ���2=NN>c�Ab���~�_i,qbRe�e"J;V��d�J���e�.�o���ުI��7S�c�h443)��r++�u��&�p�ґf�5fJ-
w��KCo�AA2���0���t,y�z��t~Mn�\��ӽ���g�E��LGW@��e��۴�	CM�Z4�����&��~i��.��4�3֦�����86�X,�=9/zC	�^��<���2U�O���i�Ğ �����IX�^��]������l���M�E�~�h����G�ZP�T�׬����L(X*H��mQr5w��J�P���\H4�7����1N����L4�\���k�F�0����:�s�W��,��k�?�f��J7�П�Td���D�0�'��^A��2����w?���n�t1x%�VѶ`V���~�ʕ�{،�TTUZ�ku��g����E_�2�Ӹ{�C*�+I}����J#��ϑ����ɇD�*a�wp�>��q;=+�6��PSU� �{��L��M�a��'6�[y�T)�.�}�%N����)��(���A�4���[zf|���໘�A��7M�$��*��:8���y�*�%���uXu�WOȻ81�%'C#�Z�m��u�����~�]�p��
.J�S,⳵�U҅<Cb2Q��������bn٣��Ɵ��:6�9i�3e�S'�CDYbM��S9S�����1���I��وG�&[�V+�B�?�����A��pgB�v�>�Gƴ�Q�BnΚ0p����E�2��I������X �1m������adG��	��i�!��~�f\Ԭ��w����g}	?~z��]�8r^q5"��S������H���+�}�)�K�g�ӯG��M�W�Y�
�L�~p�}�j�;�U���(�7�\�C`�->˾��w���ƻ�`��o�E�i[t��D���P��Q[�7ӭ�$R�T-�g"PDm��$0�Ǐ}�R|z��W,�'ф��%=�$�rZ���6�B�d�G�ezQ��n�҇�>ɚ1נ���A����x����&�3�1�ͮ�y�%���n��u�Fw͔�rt�3[GRɄ��Y?�@����ٓ0�}\�d&��j�S6:0y��/�]��6����l�;�E<DוM��s,�O��(3���v��<O�����<`��<��mv�\���f�D���,�2�]>������<'��>�gee�x?���8�D[�
�9	;ji �c�<t�B����lUJƚ�R�/����jg���͈MT�!<;g���/@�A�Ģ���<CKɕ�gz8�T�f��IP�}Mbؿa�s���|I%4��Ϧw��Կ-/ȳpGݷ�������s��x�3Kk>�LZ�Ҽ�x�r�@��^���t]J��{v���P������L�P���xX}L�VQ�c'���`�}������3�a��O�����o��'�ՑRJ~í�@L��`�!�(5�B����d(װ��%�H�Zs�ʩS�i�(zL�̲F8�6�$��^�3������LNP{�6)�\�X��P�wF����ȁ���|��d�`��H��2��7��@H����|��8nHПB�|�k���A��� �nl����o�X+�q�*��-lvy)�GJ-�
�l,�r�6�[���S���ZS�z��^!7ЪlO_�ӈ)t��A��/ʞ����_��|$�;j_�F���Րj!��k،CH�H�c�+�r���i�T��P�嫻�c}���
�>iY���Q.t�7�u|��b���#-cp�kTϠn�,������Ծ���I
@�<h����}��go�D�a���kk�d��w6����q�����6�U�+o�FWG�a�]��ۛ��b��0��[2���>	�[�T� Ŀ��?�D�k�YzMV����v�9M�����Bt�𲊊�o�y.l��9g��V��Bg����n�K�%����ӣKŽ"�#>od�����X&o��[�Ք�T�&4��X�8#����/�F\�Hiw��_Hv�>]���������dm��;:B��.����A(eE�_�Z�2���P��xQ���v9W�]Ffk�
�1ͅ3T���(R�O�]#}��n���)�k�-�w��YC\"AK����<_��m��T���xBʥ�ndH���O~d��8qt�Q7����n���[��w�u���X���e�l��zJC�W��V�de��[�=n&$�����msF�O�[-�8]'�碔:�j杍b�g/f��"�4�t�kBc&|0�Z�#NS\���3ӶN�!*�/�9%�ۅ��յ������U��u����Q�e��	����,+r�h%�Z|�L
����e��Z��_ؠ�JT�Ko}wI��7W���		�W��X�Qq��~��Bnd"���s+5�~�0AK�SO���e�!�Bc�'�����Q�#�F"�n�lo�U:Ϙ������H���?�y��q����t!lS�9
q�\N2�?�_YW��$������Z8�����[����^�A�!��~(�f�ؤ$�Ms�2�b�p5�-M�O���-h�Sud��9�-�HX�����+�f�ip���;����;���'Hz2l��ى�K�nݜ�!�3:fO-Fc W�DbZ߷��!�W�m�.{
�ʮMQ.gr����߸������G�;>�(�H��KMO�/����:w�Zg�W�����d��,`����;�ԏ-޽�?p���`�Ǽ�wGGd�c=�?G�G[���������\s��>N��sM�
�U��7S2Q�~hL����w-Ż|�'�^(�n��͢>���VnU�r�H�_0����Z���s�z��Y���HF��'��f�*!Pj��戹Q���B�<������:=��A���Mۘ��������1��Q�p�(W�d�?0)�N}Y7��3ڻh_�,�]1�w/�S�O�1�y+:񼴊�9�ش��.@�m��\*e]����m���.i��@T�}o�DUF莖Y6���vp�H�����B�f�kQ6p4K��ZD,ېm���&,g�<��}�FG���I�O�����[���;����<#t�c\����S�t��hm�:ky��^0W���H�$�ΣΎ�����@�*�������I9J��8,�V���Y(#�_��#�P��~�Qw�Wֽ�-�:�cYgh��h��Hpl���\L^y��B����n��>Ș��$��'��7�8�j't�A���zA�x^$����g6�@����i�e�I�^���q��]��ǫ:c����UI+jQ���m�t���B8�����R������z&y�Z�0�Cjd�V{g�?=��.�q�TkSX���~I�":��]�����4���lUn�v�����~��B�g�̕��5�57�Z�fF7���VTk�3�,tqK��ܸc�}��xS��>��n�}>��H{3�����J���k��Oh��]}��D�d�ݎ�<=D^����D��,�I����<9�<وQ�>U�j�\6n�I��[4����`j�t�O7�ձr�|��j������P�M���ۻ��7���I,��ׯwI��|����2�܎ưX�Kم�o55/��&�� P_�~tTқ�jl�^f_�>�>���ע����S��4~�p�uM�{�+MKP��z��0�>6����^ŷ��{O�&���ϮlQ[�ڹ��ͺ��h���{���%X����^Z�ܨ��SEc�Y����q�Vj���ՌC��/,1e�dD�˙[+U+ˌ�A�����3X���_�ZҤX7��CZo�nD>ŭNp4=��/��UE�� +o��5vr�ן��3�O|irE�nmgNj�.n�z��@��x��S�C������X��)VcΣ��k�mn�jЀi�R�]�T��+&|��h�d��������\u�B<���;�vǬ�LS�K����OhR��~%�u�����'��)���L�����OLd�Ĝ|�_\WB%(��О���.�殛'On�1�>d/~U���:�}��y���	��z���(+֔M7Kǀ���/=W{v)|f���l�&��!���g�Q�q��ɵ��w�5��h���2�0�qb�h�V;��[v���^�w�v�KS��3���	���60��=�$�O���I�w��b<�}�,k��S�L� yUv����#��� ��a/�wV�M��2�`cG:X+�_�������PF����v-��p��Ȼ�N�$N`�n��Q8�;�A������=��\������}�MCC���F��_L▨��β���E� ���!����㎎�Bk$�5��`_�kaaa����@J��ɫ�������`aU?�Z��/���IR�l�k������P��p��{�n���[Ωa������u?�\��G�Jbe���M�z(��*�˖���5��LqeB<�,��/+��٧����	�������L���8$������o��Oq,I�vFu�LB��<�ݲ�@�_e�I��a�U͑���wզ�{��S#��;�캎���>k��o�F������w}�(�>���11μ�8{���
{�e]F��7�ag��X�"ʋ��s?
����_cyn}/����N ��g�Iq�����/����5�^Bl��ޛ׭�b>�ǟ�p�p���U���dMLpQ��JA�=���C�2���U��9�>�$�ײ�ob @g�R6�n�w��,���Խu��v�:�����=#(����7��|e���
�o=���:��I���1�G�#]4cS�y���̀:����+��ѶV��*�rn��i�%�^�[ �AEW��	V��:&^]N�1���l��Xκ�FO��>�V�~�ա77K�Q�,��7���րs���G�����*����1��v��U}s�H����	u��S������RiG��j���$X��LÙ�wD9�s$�?�T�xSj�޺�	K��~�7vav�����~b#��nŌ�u��������K�!���6�׺V#9�o��e��0c�>���']�u���\{l���������B}Y�k�AS��B��F3�ޖ�\)��Ҏ݋[��i��Y�5��=-�G���'Gʯ�9�s�eB�c�FK�K?x��I[N9Z�o7T�d[y���͵*��]9h<�K!���	�?�fF~E�Tp��s�ظ��X���;U\��Sv�7�7��ه���;z(p�KSn�����<�/W�m!w�y?��J�ȼ��v�����<��0�=��������dGњBCㅫ�%=&���:<}R��$N����l0RQv��眿ˏ�^i]��R��t��^�4�]��3	�K��u��)��ąg��y����Q���X	ON�'�w�"�g�:��FWVƐ[����Xb�yQ��ҩ���j�KV��D�ڌ�΅ɭɆڙ�W��6�pZK.��ry�p[�[��*�eLT�n��np��*������µ^���?N��岒�!���%[
�����\�{yC�?��R����L���]��O�U%�Y����g6�.")�aU���m�^��K��F$�����p���������Mc"<O�ɸ��:{�9�*{��w�b�x��<�)╩�����!���(Og�<���aE��]�0JS����%oF�`��o8(Z|u��#ా��6�R�8�LMM��Y���[�mlX����['UoE�5\��=2�e3e���:1v��c�3:�����ks1IC̠�*�8�ޘP2�g�kФ���M�Ԑ��v�t�tRu8��Nlm�n������F����΢��N4#���B͵��~�!:�����f:h�2Qw��|�'������i9;�h[CI�����q��ӈl��}����M�z���H��*��u����H��brn���;�~�����+�̋(���<��4��Dy�qǎd�
��-�u�z;���'_����i%@I��p����T.E�Y_����#/|�G��+ꎫ�.zډ�N��-�-��'�#N�ǆ����}IWt᣸���*������[3ʃfd���«��iae��
t 9�|�	<���ã[��,<���.�.�5����7;�N�]"����<�N�?��V%:^�U��1a܇>�k�� cBr��3jnH����E(��]<�[�°.�J�o�Nxa�r�V�ت򆠡��߰��u��
x��[=�D�'��GGzt� ��>{���<���O8�-Ğٷ��Ϊ�yK�h�Cj��X��7;/n���(��x;L���  ).�kŬ��%[V7��͢q�@�Ѯ�R.�A���kllM��$>N֗�a�G�'��'�����������Rc�Q��)�; \[�l������zK�4�%>t�l]}U���l����5��b�=���H�t�E qg�Ýu��hc��6>ԏ>JD��o�X����8ʨ4�����[�*�D��\����\�B|ڿ+���)Gue���_��Ǘ��9���(g��d��#QW0E�@�{p���m����.e_�?�Ԯ�<̾׎	>*�c��aqy}��$vi���1
��0���V�ޝ�C��ЙO��s��]���LqIm�dۆ�UD�Tu�po�_��dF݄CY���%��{����������ki����Ķܛ�8���m��{V�3b�u�r�N�������zM��dz��$�͠��%JZ򺤅S�� \�m46lK�]���A���&�%��_\���e#�D�n���F���m�~��P�M�)�b1��������&J_���Dr�->oo1�<#.b�q� ���f�E��b�0e�8�\����;�Q*��%O�v�����aS�"o0D� j$s�/�}}B�����Y�	���_�ћ�Ï������}�D�PȐ�i�m�T}����&%4O�!B@�/�{�%�3�D�����
!��� ��0�xf�����	���J8�<�|����NA�+�ؚ��g����Ͻ�����:6�׀�mu�m�j�#�T���;_9�x�����P�-�jh�!����뒻�X�A����I#CY���]�%�B��1UJ4\Z�c���Ո8��"�$��sgy�_h�4��U�&��ϊ��|�P+�����͇\�F<�ے�?��EN�sQJu�t"d��d`�qsrОk������.}�.&�;�&�(*v;_����n�Ϡ��%!7���*3���F$�	ߏ]���29��?��B7��՟}۵�W>���������:�)��eYdy�'�G��Z�Q·������w���ƴZ])
�oݵ�Q�z�6t��oߘbۑ������O�ֿ$��l�-8�{_eo���vx|�(kM	��'�]�\0�ǍjL$%���]��T�cQ6NF����\+�w�-g�x�_r��`�fG��l��߆n�'dU&�a��ٽZciI�J���Jۂ�Ș>�]�C���t)^��sjs/��"M$�5�(Ux/ɱq\S+XELMP�n�|9m.�\����-�f�+ rw)7�z�;[Dd$tu�T�6�/��Wڇ�(��i0(X��|����/b�a�g�Ӥ�^����U�G���L:z��ç^�>���3k0����
�� ���%��F����!
M�?FЏ���+�/ɫE�ql�<��4�o� :�2n�W��H$\xX>T{���˼ǿ{`�>40����\�fD����HL��<��=�sz(���MK!�s���vaycK�f�.�据�S��
�{����hm��Hܺt��]Ϥɿa��@�(���Ӆf�Z���ǭ2n
j~�;#q�$���D�}<�{g]�"j�r?K�`�x�~8���"�\����
��bL������w�������x�L^l`����nc7��|/����>�\�܌�K/t�W���W2�x����ݬ2%P����1��&�P��˷-�cy���ê��&a��"�lO�Ѯr�m�Ye�-�HTR;̝����0�k��eC�|��҈�q��<��P��p�������a)����=�����\��5gW;��I�x��oPo{�|�U:?��I��=0��}�ECp�b��u�bɀ3�&Y���;��z�������xN���O����OpD<���P�|�9�I3+��4b���j�[��%�8#R��%�  C�,Qn*~�AvMM�RRU���^^2�u�9񎆄�	q��/j�#��EQ�o��:��SA~[��1�Tt\Z8�i�J�Ã�+jjs��Y{��c�W0�r�Z����oN�e�������h��k���/>>K��f!5*��k�`�PI������Ơ���u��C7=]o�O�C�l �B���^���lr�I%N��W,.k��kPRg�
����^O��㝈�3>X���q^�B�Ux�͘����U�>
�����h�k�z�k�Œ���S{q/�,�����a������:�1�AH�b�S���-��W�erNghNWn~ј����;�X�.;�r֐,gIr���O�Z+#`��!Vn�8م�fg2���������%e%���|oƋ;/��R&�X,�=E���r������$��<���s��{�'h�2g}<�����6 $��Oj>���:�������׆[��1�~�� �$��,ʪ���[���<���ݚR��:9�����m�'��r�8Y�HJ�ƾ�\n�q\�8�#k�Qh�֍D�.�BN�rX=E�$~��-]{�L:à8J���Nk�Ew�ID�%�0v��g��;�����J�lw!�M��#��� :�s���E�;�g�mW�5��뭜�|��kG��+s)H�+���<��:����*��p׋ڤ���h���%9�:?6A�Y�|!v��}��v��^=�����7��:@9h�Z#_��<%��Qg%��(�ԭ�*j�sP��o���o.��'8��'̷ߘ��0��e������-����V5���> *166��ge}�#,,�́���<y�9��z>�IȚ�m�9F  �J>_�M�TC�3�+��a�;[H�s@���7��e��T�r�P����/�����rU"�h^� ƭB�ؽ��簀����S�ɝ>w6�0���:�K*\o�e���>����2�	%�G0��ҍ�?t���Q&�N}����1L��Ŧ����T���ᆚ�L>����^?���2��_j��i�߫N>���/�N�x�uv�V�NA�g+��{]��� ����u7��3���t���I��&L���.��������`��/m-�a�%=�큡�8o�뵻�a���㑬�@י��&iiIh�^X���OVso44�%��M��2F^ |zrlp��"=���pJ
v[��N�t�0j��M��f�0����� �W�Ltv[�!���).�ɚ�n�	۴*��[�+"��v�1SI�L��ص�ʯ��&8-�S$���7_�6�t��Ӏ���Wy5^��\�2���*v7�/���?�h8��������byw���I�΂��v�	ֶ|̈́j���MYgb{u����U�~!%)��Y��t�y���� ��5�Ny�'݃qq���z�5P�4�4=�5	 SBئ��/��aEWF�_��i߂2tm���:7�sff�]�,|�����-cšt	X8~�����Cw?���QF8U����L��J��$����O:�-��e��4疤��У(�J���1�df��	�v0N}�,�VWp�|�ݢoi�@�iQ�8]F$��S�b���<����]�����dU)����1|�1ǤJdd�I��aУ�����M"��C��L�V��{�e�D����ƶ�Ł?�D�u# �#�w���Hۦ�û/��$��Ia�h��6}qN���+i���A���� ;=mqQC��+��~�Q.�S:��W���­n���%�1םlp�����C������q���" �齖81���/�(��Ay� �}��w�G�!QQK3��f�bͩo#��;��n�W�5na�<��l�>�{aռ^��8܌�'nXO����cN�/��w� י�h�)hc����$��Q�i�G.�1G�j����KS�]ryE���ۋ��m{h������+Jd���h���C�i}�G�ZR\��+�ܙ�+���r�9���r#0YC!&]��W˰?�K�]L8V#h4Cjˎ78��N���3�7�F��7�&M`�D�3x�&K5����O\�B|ef�|��qS{�5ccIeݙ;o�gbV�o��bŜ�3�!տ٩u�	��P'��y�ߪ���XO��;����
�<���Ӱ@��l��}����ON蠒Y9!"����4���r}���B��{%�<�Dֹ	q�����5�l����m��i�?}b�=u���ϡ16f[�艔7���1ۙ�ƙ�޺3�n�71}c��ڙp��* d3�{A�]N�w$�t��!~���=H�t@ۨx�����`Wr���{��z��8��8]����?����ȷ1s�
��V�VFk�[0<T�0I��*g�z+r2 ��I����%��4#�8N��\R�����K�Z��/D!�;f�$M�\P!!a�ЄT>�Ȃ���{Zg������z�m��ڌOO��-ʓ��*Ch�����=�[��Z�HN�'0�d1?k���F��;ߍ�ݕ�bv��SPF:�af���oYZ!@ȊJ�Y%Fά�v� ͤ�n����x���_< �kĵ�\���/�9V�Ky��o�z�����wOS������o��3�Vi�������'��������G c֬�+�sqW�к�D5��n�e݇��o9�7���\9:�������$���<�Nh��o���C�^���� o�x�݌r�Y���ַ�g��K;���s�,&i��i��L�D��=3�w�F;�ϔ]O[���>�!<f\/��'ػ���o͑tA�-��h�6��x�/[>�wvA}���ge�p'K$T)�C�,>oJY�K#a8g���h���e:o����]�����Ŕ��JT���8����H: �ڞV~ϛ�;p���n x���&G�����������"1}���Nv��Q�����kyt�4S��<c']���5nn�;�W/[df�����3��R��^���+��� �0�	(��E,qR��ٝ�pz�Ү�
pX;l��&�(s SG��� &�=�;��P�9�7�+�8���ªV_�VP0�2}ǙR��8����H����[E\*�l�l���_n�פ�A7%���㫞����g_}�]��1~�����	�� ��}�Xb!�&����NDo�����7��X����;�~��A����"^�mk��e�?�X�碌����98�By�?�b�g��1��s��v�6��a��-^rh ��>!�RF�"@�Tj\���. 6.ކ��S��a���i�@��DV���~��g/��n$��<P��y�q����}p�J�K��u�AE���VX(��"΂~1��1�yf�>HDAx���l�$Df�,*�%*Jk"��e2G���3�	5���1�����*��e�x�=�׻hD�74�ԇ�<�C��2�B�ԋ�@�]�M볁�4�In;q���t[w2 4@�(eF���>=@9^�,_�{��M߃�O���y�Ω2�C��W�s���5��~��
ķ>]�I!��	��a��D��V�t�R]%�Wh�`�'�AkD�l�#c⹻e�\NS��2�+Q�M�
wL�lB�γJX��Һ�[�)�@��R�Z�>�L]�U\F�fF(_��D�m��5�s�:u�qq�)l�5�9AR��#o�A�����tϸ������0�Ah���<̡��T�$B����/�%�煡��������'[ܰL	����	\Jy	��n+Q\�?��g]ol��[�Y)J�\�hF��d���	�g�mD'�G�{xٝ���vN��_J2�����\|0ש��ԓ�w�`ΐ��㞧�%�1�|�jm����@�_Ƹ �[��C$E{�=�57^//�R|6r�a2�ϋ+-
� ��F��	-���i����P�b;/��W��6��㹔#���:Ƀp9 ͒����0Fmf�ώ"􆈐1�̡�[n���e�5Q%��
��9�=x�e�.���IA��Ǳ܆uwK膣Ezd��a�w�l�={��YӍ��>L2�z�xl�|D��i����%,��kv�QG��t���n��J)����`��l�n8e�Ϻk�'|��ځG��|G^[Ա���L���އ��x���m4��(r�xU$��O��A���8'�ثD����k��?@҂Y_h<�!4�Ɨ]�/V�+g���>�4J���J�}�x�VPF8c���±zA��̋M��g�|d��d����~FiL��cA�j��%�@>c:�+��Fk�0{�,.�ֶi^� �(y����>p�sSx�=;;���yѿ3[+X�qo�Hql^�[o�gvGN�uM�/��f}���Is��F�*-S˟F�}�H�k{�}a��`"�d��OT����3��A�hy	O�;g��ZlS@�D��Q���;%bo�6ƞ��hg#E�U_��F�A�tH7�)
H)�).H��(]��t�t#���� -Ͳ�t.������;�2���>���|��y^N�:>�?�+�mi�|��eA>TߠT��~0??�̟�o�~�	��~�>�������d�;]���W=���w����Vɳ�zKs�_�F�,~"`S��u�kRA����4�5>���%	��_���~b9�+0_u4�:8�h!w\������c�졏��'�e]L?K\��5���vN[<�u��H���ʍ���{�gU�L���b�PD�#V�	�9j1�F�|���qv̛���u˪��Of��fQ-Q3�)����QJ�T�5�t�lR�]D�`qÝ_�Vۗ�O���,n��X4���u���	h���O&	:e����JZ�$al�}g�H�#iQ��@��3I�����F���&�7�lFq�	g�5j�Ky��1�&�z"����
Oz��^(x8�%� ����+�M���%lm�}��N��w�ҍtw����r�C�/�q��̖��Gs���`G�k�u�!)�V�z4�����j�%��+�д��f��/���j��K��w�����nj�l���ߴ�����+�W�x���2/�p�r|�=a�b��'��g�����*������d����o*�d���x����f�ec�
`0F@���]�_cZ�i����=<���$�	��>l+}����7}�u�퓍�U��(�.�OO؞����0ER/�`�0^G��,���Oz=!o�X1��r�z�g	��ڊ\�����*k��K/K���/�g8�����{�./O��O��`n�&M�ۃ�+W��ʬI����B�0� n��+�
ד�F���ʌ	*�~��3O�/�G�J	�1X�-�����A��nͼc�zXF�i�7�C2�/e�6���N���#�6ǸfS&�_9K2*���9��PU� ����pA	��oO��
�6wB7��xK���3�TjĊ#��0y�H#*�[����.�V��v]�x�>r�Ű�w,L%���G������*wh�QĜ��i`vl�ߛg�k$�=	o{�֝��eo&=�.�g&�Ұ�l�lﷵ(/���4��+O�0l�Rݥ��`��$S�V�<�LtҁtWJ!�f�9�o�������bf�u�&��kjK뉢�̡L/Z���0;��L��������+שmwZ�2���4xl�;)�8{e�'j ��ۣ�M���:=�.T�Ѐ��H��0�.��������1ܗ�L��ó�?�/�F;׍��J�iᗕ͠�M�
��-��J��	 � ��1J����ܢ��NJ%Ծ��4M��`!�>�>⨞u~қ�)��S���V@tt����:��'%%7촋F׷�F���}Q~@W��٠�lXǏ�A�Ȝ��j.�Q�'��y�����'%%a`t)���	RNz�1���?n�>��*v��b>��� �/��1������K���l���p}���r�MҪ��؛�-{�9�R��S��﬎��Xzׯ_�5]rH$r\��֜Q���v"--��2�Z���}P+n�&�=�U�bV�}ʫ��yN�7��zh3�O
�Z.�:��̗�Gmٔ=�D��o\c����3�4���18��;����o��?�`��>�>���B�s�(�]����ǃHܦN]$��R���	�!Ѓ�RD�G�/q5k��z�$�L��zj�3�5�t�%**ՠ�}�ֱ��8"˞�c�Joo���`8]r�E�� �v�e,t3B�sn���\Џfu��ҨX��9�0��>=q�Oc��7��/�(��j?r�������I`� 3L
��Sϱzܵ�>n�
 ���'ω~h�9K����$��yм���U�e^s	����,�b��u�+�G�Rn�<A�m+�F�V�3R2�9D�:��̇�������桁�\�G=#��R^jglKn���w`խ���+����w�^[y|�(�SU����������6�����+���er����7�.�&�m4�wu�5M�^� v�I�((��}�ޣ\���=n�)���-�L#�h�dۋG?\����4�4O������
�	�*s|Q����9��J��~:��^��ߟ�Z���$G�G��]��Z�.3�E�_`����O���,�PN$=��,��4P��y��u�K�~�;(�|m2��|!qT�!_	�gy{7�� �^:�1{`�J7!:��'��\T�zA��İ�����/�N��*�j!�&��xG栗RP��=�=#�aΣ�W	J�۫NT���Y�z���hr'/It�J���T�{����u��@j|�;��N��b��S��?�ң�?8��f0g��t���%�d�s�$*����ћU���B���٭��?����5���uӼ��ʀ��r���W�Ύ#9&��ݗ��]�ß(Te���^���qG�E`T�Ys�Ik�Pgp���B�L�rt`z�g�h༖������ך����3Skf�ד+�g�M:rHZ���l��'sxyw�5��< �d�&br��/���x�߈S��Ⱥ��Q�g����JK��CV�V��)��e�u*�҅�02�a�[0����c�n��hz�|(��@�9�/��^X0=��%���x������.a����m��UQ��&0��?�[�yy��� ����	fMϵ�ټ��<ݩ����]8�Z����������fD#���I؁�ɺ���8+nӆ7�X����α z����D��yL����L���ͪ��S���� ��������(2NAQ��#_,���Z1=e%��;�QPS�ۯo�@֤^���Sֆ�&l�(�+�O����hf�W1t�J�������SW��-�]����_4Н�a������"��/�;;Y�C��4��0CTf�-���-%��L����ϊ�`�.���I���G򀿖N�>V��gK&����4mx�x�j���.��5p�J�^�)帯�A�1Pm�?�	��QjP�֫���ο1�4x���|�?�d��&�V��cA�M�IR������)����f��ͫWM.	/)�<znӭH�uuuj��[x�����OA�WC���˽_ ���lf�bIX<�_~��
��������t�)�b�T7��ñG>�{~s7}�1��b����W(�+˿["8Iq��h���	j����n�����@M�/��c��9�*"}�/��jS~P�8�{���r��o��
�K��^���ٞv�K�Z�׎���(�����	$�ڟ��6�_$������	8��TZ�d��z,6Y蘿��	�#������kX�BЗ@��g����=_�0˩�p�KJB"y�/����D| �f���u�sj���t��s)�7��U(:�֪֡f��ww���M��l��?���U�>��R=�~x�zG��W��~�d�e�ե���s���6���y��p���d\=QB�_B�d#�L��3��]2m&�i;~��2Iqѭ˴�D$$p�����i�&UC3���.6��Z�!�હ���+�v~�X��o���O�N �P��K����$��&S�ne��25/�v�$�q��az��ʾ�d8eU /�iT<��bmt�%H�M�����Ә�p%oP���k�|�8���m����qS�4H��^��bLb�2��Tط�nX����?�u���z\�Pe��U�<�Ү}��DZ���C?v�*!��4̢t~j���E��O�?���2tG�F?f�T�avW&��\%��B6q_W�L_���B�ޢ���ۈo�vj��X���2
�u�x��g��ҵ�ǷL�C�sS������q����8��|	.�mX���}�D�u��Y���mʃ�K��[2�d��>���;z�J�����?7;�%�htf��y�j%����=Ce����E�0ڳ�clek|��J��b#�m��ҹ�����A��]��C�[��sD7��j��;�)H��^oMb�����Z��w�U�x��Ȅ�fP@`1;�L}��mp7�A�����:Qx�9~��i�8tvLH�˔���t�P�� ��)���Y�㍝�S��ț�N"Moӛw���ulm�"��>k�x��AgOlpr����I�;��u}�w!\*c���.�(~SV)1�����������t�O�V�a���`��8�����,9�+����z����sA"}K�n<pd}?���Rz��!�&�t���b������So�ĢP~���ë>$c��M[�R����=���k��'���G�`�bg�����\i����B���Dڂyn�R��2K�Ϗ��Vwn�����2b�a+�`uˮ�o�$H��������ӾR�ܱ�D���$��%��G<�R�fj-���X�-�RJm�H��{��8��XI�$qj)9�A�/�~+�(y\2Be��=��@�5O��J���/�9$wq`�{�-����^���0�vzv6�{{��+�I�[�rE	�y�s�Z�G7�z�$�[CXgwQ)��C�b���B�����P�u�%Fq�Ge����)��usV|�eCRB-n
Ov�ަ#���y'O�}��	]v����%a;CD>�S��[��3�RN�!	$�:����XR5�\vI\�t�/��*��A]��<��}��Ŭݞe@���_Cg��l����]m���Z��YA2�9:hZ�$g��R�47��5��(.�@�XtJ
~��m.���s龺ݹ��$5���\J�1�Ҽ#`����n�K�V�Mq"�X<�V�9�8��n��/D��6r?��J��gV8޶�V�T�z������"[lf,�'G�����U�����Խ%jo0k��@��hM�"��Na3��s�o�x����a���1�&�vv.05;{�	o��q�r���Xս�7aByF�\�W/�Z��vv�|�C�(K��ڸGts����Z����0�c����as�}]0g����	�{�@��KM��l���lr�1rx����6��e�r�JL.Ԯ!�PBϩUpxTi�?����_�*B1��_"^���~�2��fO� ��h�~�.�����8�쵺=���V�K�6Oe�%�e���(I�#���t�t�!)��"@W��oN�6��Do�/��J��o�B�,��W��gBKʘ2�Y��<O���/�̓�����Ѭ��� �_[�k|ef��;�o� E��]o��2r���^����y�߁z����kh�~W�}�LwG�݋ɞ�M����^D�9�M����k�_����~Ҏ#+w6�(1ѿ�]����+��d���Q��L�X<��Um�/
w[4(��CR�t�@L���f�.|o��VO�A�6K�IG%\���Df������ck��)_*����4�{���k?���j��NrЏC�%�o:��(�xH}��fX�:��I]�Z���sN޾�:�����������o�LDtW���r���;e控\�wk��X���l���w��l�����$-����v�;�J�BW��!4���H�S5��s~/���vg-(�^eċF@I�6�NfȞ�l�>�>�kd��9����z)�������JEOO�{C�y��ig�6¼���rglt�I�ުZ��n]E:\�3�<�j���6�s��W���I��M�qK�"����e90����W����c\LD��g}���H��=�`O���o����)f���96v�S�ۅ��%�>$��-~�?-5��1��E�$��ޡ�&�8��9���ou2<��U�lݔiH�����cz�=	�K���c���'��d'E�F+�WM7�0*iկt�I�[T3C*��~�	p1���s��v'�_�|�u�:�Y���u�B��T��T�k}���Q�O��:s�����
r��w��)�wf"�^E!�C|�&��B�J� .��.�}\X���tB1�៙��f��W�L��U���*wPki=*�3���q�i��)�rN`m"��3�$^3��X�d�����o��n���<�����x��,h>t���� MT`�W���0%gp|���Ԓ!F��}�ao� Z�^!�Zx�p��-�fM�U�E#(�����˦`����&)��沌�K4�h�,{~d�ϫGߍ������K�m�^NVA3>����D-����Sծ����'y���������([��88h3�h��`@lH�o�k�P�шG�@U�y���k2���U�D �lȓл3��,�!���������ZR�E�-z1�_NT��؎��De���,5�$�����z:�g�z8����į����G��j�'�tuu#�8B��p4G�f1m��ނb5oW���s:Sc�Fm�|�D��эT��^N�Laʣ��H�x��є7�u>eh`�j4� !T񋋨ܢ��%�������C_���)���jC�+�J��z��bk���H$>�wû�➸,Z�x���K.�lV��D�� j���W�BE�6~�e���Ncͧ���Ks8xj"�KՈ�w52�
x�&6���yl�P���ow^�I%X�#�h��ݨ��W�B?�͘m���pOPH��+6�����L�7��[n�Td��)��C�௦���3:���/}�Ĥ�^��!���,7�譀�E�e�#g�̯I���.���S��6���5�c�<K$��0mI9#u�����?C�ȶ�٣�B� �m�����\���Ob�wIȊ���L��+(�dw߱���1���ߝ������0�r�n/{N`��s��r�~afV!E|%0P�L���+�o+$���I}4�mv��9\�J5~jB�vk��q��;�?X���ᩒ9/�ð~H�7�((�6�6w�����W�'�s��	���Iț�?�7�B�T��8���o	}7yҏ�_�qR3 ފ��poC����sΤ1��E�x���8%d��T�Q�[B߈��tW��8e���	]����iS�I�� �Sv��U�Y�$��5��0?T�
I����^��UA��^B���K��׸��R��c��K46��Kw��4��`�+�
��'����튍�8���t��N�4Se{�0���&�^����8�ק\��EBe��0�����,��!����
Ǝ��\B!���&�!�X�4�zw���>�|��3ڬJ��H�-s���g�/���=��}Z1������|Qbb�]�k����ڡ��|���N#��+wr?�
�i�����`��$x@��!�mEg���1�,Q��f�1�dswY��.�an�'\�;b�,Sh�dG5FPL��v���0 ��H	WVV�Z���[5�p�L,L���Q\�'=YIH�����wk�kD�n�<����L�j���C�.ںl���ġ�UvP�Xp�s ˩���qB?��� Ōf���`����6��^S�oꪒ������h�P�\�鿼���;���f��
�s�����}���y�PyѪ�.y�������N�i�+�Mxk��w�<߯j3C<]<��O�p� ���A=��<��ތ12�(���W!����h<d��Ӽ��.�̭�g�?�Hgc҂�ؙ����d垝��K�sʬ����)�rf6!M?/��3|�g�w<쩤�"1Y�̨�!�������@P�ʱ�$��}das�2���Wפ�w�M?E˿ҿ�a:�4�ů�/��L,�����G+�-7�@/�~2�ؒS>�Ǧ������;c�=��Lݓ�. ��"�ܦh�J�A�d}-͔�ʔ�k�yF_�l��DRٺ�G�3������1#vc�� �8��^�6=��8m�.A
�4oY9-����q�_���l~��:���k�� �1�_i�|�/.���"��Ռ�?�c�}���p������_O�x����!�6K��5wqQ�5��<���/)���2$%L+��������ء���L���RM�޸��g)����?>zA����������r��m��KL�c�&<��s)`݆���.��r���6mI	5i�D��4�_���o��x	�bO��ʯ�av��T �	?`�c�?�$K����KD�ۇ�a=���yRm9�7�i,���n��oO7�j��Y-gH�o)K��D&�q����#P�f�?��L���Q����C���}�7��$\��ր�ш���S���,���J��oʸ$�g3�ŏeԌ���}��Ny�����/h�HiU]ޥ�W�Na���`պ��o�3�2���]l�/�6"���V��D����o��z�����Ï'��<�)4l�
n��{H���Ҳ�+nm�^I�?����<>R���}N �
xǧ]e{'в�U�z��ן)M���+kt*�
#�5����� I# *��:�L�m��#��(����)jH��z܆R12�D�-��y Udx�cI�� ���6ZA7�s��\����/�!�p�=Mf+�9h0[2��-��u8�y �AbT>G����Fx!(㾡ߠ�`#`��[�)1�p���̦���-o�ct§`O��YT`��GTM��C棞|�򋷵�0pQ*`t&�65�T�w��I����9��B�����I
=U�;6x3O)�v�����cD&���כ�ұ���5���r�z��l7��s/3�r�J��0�<������������"TC�"'�p6�f����(z�q��m�N�;�-���/�a��W�����I��t�pf�HQh'��*�2��%���"f���;���������q��J�	`,WJG#����RO"s4���"�/H��Yl���8�������("�KbY�{�ۛi����a�����]�|ӆ���ndd��~'�!��D�ˌU[��ޔ�8���8��Z64d]���fH��S�D�����J1P$�`u��5��H ��F" RS9���IQ��.�Q�砬�2�:B��-�ȃ�s���ܾ�K���T��x���+Aw6᲍ݭΘ�!@Ʒ����"Z�}�rM�@�]Z��Y2h���٩A���O<���!�S�d�Ƕ4y��##8g���<j~�f7S������C���5X�Ϟ�Ȳ�ʝ�g ��&w�����N�5�X���lܯv��X0��M��-9�}yԫ���&ɦ���T&Џ���x�î6�	��hۼz��\��T�#"�xҭK���M�gI��p�Ͽ��9��Q++��B!�"��M���|�b��h�*O�J��f��ު}}u��Y�@�M�!##P��]�b@�um���O���DT�FKG��*�VH��|�L�=�نm),:�5l�E.�L�7!��v�������vM�ߩ�c�S@ޜ���-,:�MQ"B$���@�jo����DG� C}��Ϟ=s��.Y�t�ś��ݑ���e��;�O�x~���K��y�x��~"�30�k�e�[�$���(�_�--M*�pH�����e烏7 6�����,v9G\�{H
tJJ�D`�"�W�ؙ����Եy$�;�&=���B���A1���CNa[��"�s��u��}l��2�,�C߻<ȁ�����|�s�>���B�_Bߛ��W�BNr{��Kn��v�zV��`�@�$Ӟ|���90�j�&��F9x�[�D
'I�S��|RS~��N�;p�>kǳ���fj�����lѧy��vl���
��q�G��|m����ǂ��̬%�t0o���۸P�<������p���MyQ�p�^��V��M����pKy��'M1��A��������صq�٘���Om�ޚ���?��b%K��ӆ�U+�d��O���Y������Ŧb3D��L�����FT�3W)���̮o<��c�
���|�K�lh�`����FF���|��26��L˛���'�$P���CRrZ���5�<$��l����^
� >j������
�@FMV�������f##����oU}�?c��˪w��о�A�s鐮4�����BI����F@+��T�z	1Q�>�U��o���z֒����Q߬�iC6�m��(NvT�� ��U����ɴ9�����H�k��W�I��^���8,��m��}X0��F�MNB� &=-�����d�󬏪�yϛ�5����������
NQg��ɰja�`���:��f��,f�̀!�Q�-�q)�'fJ�4o��	�-[���Yb�O �T}o/ i���Ч2���ÞH ��^�o�f5��� ^B̩dҧ�w�^Ǯ��������
��`���!B_B����.x?_��Ĺ��_�'i�_�����Ʃ
v?��]����������q�o3|H��P��2$�|��[kl�iQ9�,�������&J�@U��w̌�Nn��un�-����[<�����x��^'8�����I6��"��V������`6$��0�������G����U��3Q��x&�}B����ǂ�� JbXV=)�i�/F�[��8��7#�cF[e�==@iՁ����u�/z��M�6�PH C�C��p��~{�g�n�`C*�s���$5����͕�`��T�M�wm��Kv���)B��٦ |�$ގŮ�"�S��N&[�:�?_驺g���H��
rssf�YL�ͧhYA&{��+aǊ7�������e��-? ���M!����"�r{f��A�������r�	�"���6CZW�o�7f�!�Owf�)/hz�gQ(�r��{;	@����}Q��8�)-+C �5�*��z��iK E~>(8R�r��3�'����|��M�6�T@���1m2���R��.Z^"*����N��IT���y
*e�\����K2�u������/�4�*�����j|�}M��n��6��Y1T
ȯFR��	~y�a�x+��裢/��biUl?�E��������)�uo[�����Gm"�˟M��O,VV��;z�؏�b?���&�l��^�'
�'{\>�6�f�H8��&�}������F$-�,�	ȏ�����]�S��;�Q�,�.����� bLj�&�۽���L���1"���T���2��0���.���TS���s
��;8���sC��4G]���L�[����ҭ%?�խ�ݩ�h`(
��w>�f��	��TÓ��[ǭ���'{��8��dP�55��C���<���� ����U�Rs¬�ͻ��/FEBI�r�_����P�~�H[#�*&�y��^�{H��6 ~{�{�%�s:V
xN.���߭�X-g�醍N��iܪ�g�T㕁�;��h��xG ��[�UW.}H���߁ر�IϳۢӾ�������ls���V������"�Ņ;&�+OƏZ�o�I/��<�ř��G�r�j)�S�GP~��d��~f֋߂�~c� x|~yy?=�ݭ���-,(�����	�3�2���KVD���.J�����Ӓ����V�l�;�H��1�Y"
+��Yj��OX���uu�B���b�t�����!ֿ[/��Ҟղ=�'�3�>9�0�$�pf�P~_u�T�����񛚇c�N����9��<mQ}��1E�&�V���uboM��gk�-*kg����MQ�� x\sPfq%��ۦg�,L`f�V$g�&�ܴ$��cg�KcQ辪ݒ�C�����}��<�0M�@����v�F�-W&��sc�A�M�����vo���4�@�S"���ʝ�����۟Ar k�2�`?%��.����Y\f�mDLazd~�َ�w��hF���F<�]�)�O͡������Q�Qp�Ic��wnY�w�W#���gC~ȟb$������4݄�0=T2��f��:gb]�h���_h�/yJx�1}�ʹV�(\��7i׾���ѥ����/-/))iW1[*)�4:���Sĵ��ig���N⓸����������}��G&"�+s(Sq��:���`�����]5q,֥���B�i+ݟ�~���)�߮�M"�koW�t��dsT�KF �	�lc���w�"A�����ˏ1��}�Ɇ��z�-��h�!�Ϗ�"���y����A��H�ڏ&gC������F�v�n/�5��W�69.�ǯ�oQY�.B�[q\?�P+d6�)굿����-�;���v��bs1���'X��-�<�,v�������)�g�Y�H�Q����4�B����蝧���6=��O���}��?�O~�a2�WPX&��'C^�S�b����VU�ʏ�+�"yg������2�K�Yg�z
:aP�"����_m?ا2b�r�'(�R���*�f�r'�f>[HPP�X�Ր�����qR�������r��J�Np  �O�#�B2�AQC�S�����P�ϖ[��s��URҜ&x>���}b�gsl�'r�7�y�Ec�IM4*wt����p���kE�G����"y��\B۹60?XK'��t�H�����ة��B,"���	�^�dcB۴U�Gh�+Iw����,������g���l4���a���MQU��-���Q��f�_�~�)�0�䵴�]<؆�g�ZRߎPK��Þf�4u ���Y�\z t��(�g����c	�91e;�x8j����ڭ���.?`[\�(=J��rRy ��q�^j��F*Δ�@J$��rՙ�+�
�Z��ׂ(ORH���-q��+��w:�l�D���D�~���층���0�`]�J�i�VG6�Y�Q�}#[ku��FR���wT|yy�e���A���=>��=tc���[-����~����˦�"5�����G����T��)ξ~~�W�*�ff����aJ+6�����:%�:%_?��z����=oiKPT�M�����o��XN�˓�A5<�u�Jj����E���,''7���}��}f!y��Ԟ���K�'�O23��1��?\�/���Zj��kp�ڥ�b��r�PJ/���p���ۗ,����#	=�f��d����^���!�����-S��j���O�@����>����s9��%�kF֚�f�L����[�d�PlE(���v=t���B� �����i{��s�0�zEG<郮V�Ov�#�Z�6%�פ�7Cm���1��
�ϩ�?0��/3��T�n��=U��>y'-d׼Y�*Ruj*�A������cM�����b�WɈ�( �$T56q��&'�/d���c
W�uzcO��Ч�K���Upb�ׯL�ϹȠw,,���\�5֐Xܠh�&Ƨg�В#�77�D&�9����_ۯ�
���1�{^���e�T�B�o,C���빼�#]Mc����D��"EϮ�~�6�vXPN��
� �����OGp<�����*X���(�r�\��,��¨�s_�����R����k땯���ŗ�KKK�����U��V�����C�M�66�w�?�u���z<�e�{�-b�w��G�uuq����匎��g+Lͼg7��I���A�%�1��	b����2q^n���T.��R3���K�-ǎ�����L]ZZ��:��?���=$@s��!�pe��kcG�]D?���1���6��9�˝��������I����ЫgILc�h=�A�>����1n� ���h˵g_qZf���/��F<��M�>*Z��eq�3)`ڝ�M�@���ƹ����:���;��|?���[R��Å�e�����,x-N���'��k��Q�M;�i�gҧ�>a�HABB�����]�Ԕ�뗠�guC)J�;?�X	G���/ܜ�<��d�+��:Y�R�z�6����p��������4E:%\��x��  f��s�gk��;z� C�*#.��/�]Er1kBi��!�o�&��[���ʅ�I�k�Z�x�̃a~��	���a�2�d�,�Mj�b7�����d�@��O	�����e �F"���V1\��=N��o�bz�E�/�J��{��D$ͧ;ס�/�Q*ϞˋF:î�n�.�b��c���*�������/΋�D�T�%.�uי�[^� \�w�4�q�+/�i���`f��/�49��Na�D�!5��b�&<���,�mHe~m)̀��ڿ�½3����'�wƖe {e˅��ݹ�G�FMԀ�{�7��	ikV��*G���j���b���SE8��e�>�A�uK��5�4Z>m{HϠ ��4�Wċ�5����	9�J�`+�����P��B=�0867���N�[�P�^�
vo��3f�L�5]%i��)���m>^HT4��p����47w��@��C5^?P�^��ş㶢:|c�3�O'M²[?-���g��o}}}	ZE��9��NP�dSII	�Q:�ysl�p�h�H����$����BM05(J�FT�319L�"��Q��>^U:���	N֐q�0e��ƚ�6�E��K/�:�a�xF��@R���3̝��a�X���H��'����L�s�=��⦸IE51)�.��p���ƷC����<��q�E+�eJ+���p�}y i��=�M�.��uN�3�9�r9?�?��rT��SЩU�"Z頳(;�F�*\�j��<߸�=���q�|w~�G~s��8��5ݿs��1Y��㞄dǑ]�6i8M�E�?��2��ňw��v�4�9�S�9�>���)H j+�"�GMO��Y�0�`�h����~�^;ȏ�ZWz��M�Ǿ�Lj�^��(뾤��Ѭ��*G��	�L����m��#t������+Td���Y�Y8�8V��ER�`lQI�4�g�7��!6C�f�o�j@�Xח���
���W��b��XϓO�`G0�b�t�a��e�.DMٳAĜr�+++�'�8�
����O�%�h N�:�F�?IO�%OP�b��j�
ʪ�x?;*���I�j��� ��W�D2���Kdzy4���!�)��IŬq���1�r���� kq���,f�љp���u{۟)Y>����oB����{B��^��[ �A�w��v==�o���ill��*���H-�W�@���8[� �]���F&�r������#�2�+<�S��_�4�Fv���4`�6�t
�j!��9���#�{��_��+a��.��X.�~ᴸ*�������3ҩ�e�pi��=�,�x��B��ژA�ej��2N�_i�(��R��M��1P��㸉��r�=�r��� ���ݮgn�M�YJY�6*d�mK��[��'���;Y��4?�����<��LK:�s@g��il('?�*.¦���6���7kw�BJ��Y�����݆͔gw44�M�0�&R?55�>���p��6�dQP=��e�g��%�&E&7WCX__���O�%UU��L�΍/�FZ�*���?�����W�@�g��t0�ǭϷG�x"��l��.+ߘ��G�ES��(�;ȝ^<����LO���'*�~�Y[����%x<kb���ic�՗��c�fy:dmL�.��)��x�b͕�߿���o��:~�B�z��3��%�_0�'(D��)�
6b<u�Zm�)��,ە��nk[/�9�c�[4��E��i��JOX������s���5���ڤ�4�Q��� � |X\�no!1�s^�C�w���'-�C��k�>�l������pձ��m��R��~b`<����Xud͵��W�i0���L��5Ng����5�E=?�h�V�5�ޱC��W/�,�~7��$�U~\ss>��$QO�|1*�x��2�JD�J2����]�XW���}�͔�'dz���Q��g�Ⓠ���]�fл+JyK���N�&�c�b{?s��\L����w�s�^H��I���p�T��������V�~(��խM���s�4����m�`�y-���P������^#�[/��m �%矁�=2l�lp���'-y�x���w���]/�Fm��w�% ,N�;�Ⱥ�ե�'>����>�=�z���߶�xk]������s�����(K#�H�Ji/uj&u��]�P�dEW0&�ߙ��B�pz'��|7���?��U%Z!:��Ѭ*q�:ؽ/J03�_"��
Z��Y�2��<iA��)&��ڛ��iO����o�,R�q�t�cv"X'��ɴP�py�����I{��g5U/�elT�2<�b2��������0��ppC���v�t4+«���LsG�FU�.�A��q��*kj>���M����3 �F��#ej/TU�[=���z��e�N%���G������RS�DZ g�7a��{!|��p�R�޺�	� ƽi����1���}{[��&�$���pJ��B���C2FG�M�F\��.<��6�rlR�P����\ �����6-�~��VQ�'��O��&�0�,R��Y$�.� ��Q�����	|Y�Ђ5/�x�YB#,���q�MD��Gإ5�t�+}���P���i�������ƕ�uz ��q)
�o{���5�c��qf�n�TgQ�4k+� ��׍��Я"�w�ъ�[�iŤmt��ۅ��B����	tQ�y��!��g� N�U��EY׈� 4qȩ�_�Q��;�ׯ��y���'��ǫ�X�Ť�]�p�;��K&I�;N��ޮ��ωK��o߅�H̶�9��ɛ�F���D�oW]^�O��TEj��,C�?	֌��z�t{��F^6@u��b�jH�H�-���~�pK
����
=6&r{,&�i�X��tꦌ��5l[�,�U�9������v�, �l��K�B;ś1�u�l���MgVzU��W�"x�o����Svе��,�����ͽ�{��&p����2U�C���XO��A�������چQBR��Q��NA�Aah��SJ�N钆A:��.)��n���������pf]�>c���M�5�*Ua�~�p��2#�wJ6��1��,:1�$����
����j�i�}ϣ�A{�n8!��x�J�ۿC���)�CTXXX�v(QktD����腩l~�}�����d�d�Q�:���U
��?���\��e��74��kqc���DFm��a�~��A��",�
P�b�p����/,��k
��\��ٮ- ˲��|�.���2��sV9��|�(�Ӌz�nd�Z�ۤO�c#}/��'���^������f"m���hd��V��s C�}C���sD��)�$<�=�>l�7��(�1~�8~�ȝ��\���ƀˠ�ͫ?q������S�z� tt�!B��2���&Y��Z�������z������G�#F�E,�3n�xe)�w�Yۄ �)��]�B
(LC�����L����I��e��F�+�'�xiv����OmZ��C]����`�v�G�\_v��a�y)��{~O��H�	F^��KS���/]G�l3ª M��%�^���ῥ�n_�Ev���pw�?T���N1�2HǨWR�gv��z�A2��W�bM�$j�~����n��n>�b]�`�a@~��`o���l^ e|a�?D ��Y��1�`��N�8�n� �o��/1v>�Q��.� �>�_�?D�rQ��H;�cK���i*x��G�C�O��7$����j�����6
��(?��\ ���bo�&+"� lD�G��\���֣f��;Q�N��v+H��ijc���$��K��S<;D�>V�����R^�Ƥ ���5��(�p	�����(��ܕS����,6}k������?1%�9��j:�t`2��h���!×��:vuۚ�E��Nc^#q��P����Q#����;��B�_}cn.B��V}��A�
�%�77�l��Ǒ��|��.߾���"����������>-�ã:}�#��x����HrWG�B322�N@	�^�H�\.9��\I�^%~	�0-T�(l����d����8�?�KlőD���[��d��ϼ� ��������Y]�}6���O���D��u3i�`_�j�vM�?)�HHͣ5ƿ�,+32(���3p_��ӊ��V�O�%�+����ܡ������ I^	�(@+�%�;K�K#~�}����9Gʧ\�b5������-eaX��^J�wP���9�鮀=ےW����S��~q�/���킼�CAV�^w$����Mwg\�:��g����'�i�]}��#?m�s��']�N^:Bۘ�5.�w=�7�� U��X�������"|�QbW�.�׼���wp��4<<�1����I���&�
?7�"����U"�U�t��́�p|bj:T��A<)Sx�Y��c/�4��Y�.]屫Ӹ㵐��G�X�s�]5��'�`����wz��},��n�|)#D#��J�%�ġ�X���������>R�W�N�Y^!ۭ�U�b�z��H*��s}�O��i��[^����k����s2r����p���*U6d�����g��ݎ�_�W;6̴,�J��h�zNj��y���&>����`�u���!wiZ����f�߳1�i��اy�\��4����))K�����:	�K���kR.�@�>�����js���K>����x�JD�"���R�����M"����!u!�����^� #�����l��2���Kp�Q��mX��;)��xn{:�����Z�%W�B�	<�����}��?�1<O뚂�bk�&p�@���/��eCJ#�]*��<�A��p�P���Р�!��ɰŕY��M*K0�W"��7#c2:�l��ڬ�6�}C�OX���^�.'��ه\��5:��CbJ9)L*|}}b��h�C���j�N�R,����y�^���e��ʆ�c��k�9�X	 M|g��
nu���y�����A�?l�Q�^��\Y2u������=6��ʑXܑE������vw}3[G���U���\�ZR\�9�j��Ď��_����`v�do�h�NV��:P\\R�Yri��~�V8,�Xh�7H�T/�w���د��(l)a�h�Q�s!:k�-�fe�A��yV��
�B�))����9� s���H&Qթ��3M��g�B��/�R���Xt������!�j�d"��	�N2S|b{<����&{c\j*3���ij8@���	�A��TP��r��$���Ez7w�N��+�6�9+�TP�7`�x���ޅ�U�#uvv6�R��U�^���ڲ�aV���q�������O�L�
����&����Y��;dz�����O�(&��Imgn��Nt�C	q;Ġ���xmt;70�ۖ�D|�)�|�d+�;��c�75mk����[[X	���с<in|!S�k��;{�}�|k��h�aq��\�PrU����Q#BG3��3Mʞ�"2p�J�j��L�%OS�uJ�c����vb�E}8�:����4G��22н�I8i7���R�57GS-V퇅�C5����+�Lcޝ1���jG������海Eb�^���|��(�*�Qu��E?+c���y�u>Ͱ���ߐ�ޒv��sVF��E);�v��*���.���p>H^7l����t/+!zD�G�l}���Q�2>
��a�cz�oKf�-���N޶��׽j���.��z�����a����m�or�\��LyB�VP!��ۿnF%Ir�/�����;���C2%.���\s�ejCq�޳9�j�3����-��B8;`y/�>��6�M�T���������蠹{I�+}����J�CԊd::�KS�,r�WQm��lgY�k�;h(7\�}�ޏ*�3j�M���8�8���$�i���,:j��Y;<j�2K�KB�"?8��xHR.�,�(���yO,�h�+�����g=}*E��\�rA �	���_j/�Ş����QS�j�5b�]���4��/}7��>V�p_s��D���2��4�@}!I|� �Q#ǱUR��_]g��=�E�&.�v��$�=�׷�������.�il|e��y	�b.����u�D�N��9��x�6vϯ�4���rrr�RR��N��c��T༛@>��0?S�>܈'�)���p���V��̜5���:��켏K��
�"mU�Ǒs�avz��f���=��=?�낣W���6$�E�孛ە�K�ҳ&�N��z�\�&�.�:���}��T��)��-�iN����#�|A����k�N+Z��3���ǰ���;.S���G�8��$����q�6<��L�[����p�t2�>��|rQQ�S77�)g����T��c����4K�ٔP�	4��4L�as�+#�@�К���r+����7�D| 5����6]�r�SZ��)�M�l<=u���68��6ihZ���[�:x�O��ZB.a>�Ɍ!x�ū�UF�?�Wχ+Y�z|q'.�u<(z�्MJJ*�v)�n[辤�xȬVX002��ly5�w�u �,j���'ʴ��I���� ��_<��^��&�sY8&�K6�S
����ċ���l��I8m-�$*�n�!�@��-���
L�����"�_�fM������P���.�/��D�AP�E8�);e���!D��5�9�n����7�Qÿ��F��8A��\w��k��Ri��#����Ś��)[�B�T+Q\&Sab+壼��e��ι�n���w�B���v��s�ۿv+}����?Џ@,�WF��}3�b<��ϛlq����6��8��g�$��Qj�h2r��Q�Y�P!�BXճ" j%�XG��8*�� r�̂[���j8����}��W��P�{�P��ޖ2`�A�7��L<�o���I�,��w�aN7a�v�7�˝=g���(Uݶ�����y=ޤ�7h(y�MF�$�Fx�Q7�z0q�Cq$��5�w�&��4<�J������]�b��3�#�]i�ۡ���Ն�G�/`������(��3Ieī���<���^��q��h�\ӭ��/���+����_{}��2��)��}C��E��ݍ��0_Z�a�4��y�\Y�X����L�N�UTT����V�'rx�Ƽ�O��!u�	�<�
B%Ǘ���>�kǒzt�� ʧ��IbX;`NZ �ą��MɅ{����2-�GU��g>��ʒ#�(�]Y}�.����L�%$sPS
�|p�ԐD� �M�e���/���ĂJⳀ;S'�>�9�� �P��}���ǵsm� 'ܕ/�+%��3�+۔41jy�O-�7$e�N����y���%�E�S�g���C�	�����@3tA�}��͍6͞�|����A�~$F���(:T�d�e�L|��M����	m��i�^��?��ݹSGQ�!S��g3�:������X���.hO�o�p�[c1سu����WL\�8Yʢ���b�?�	ND�Ql>�:jX��
q��?���%����#�W)���W^�i�w�P�WZ
�d�5���J|�ŭ�QB�� .~8	���A���6��D�M�Zc�ޔ�Lx�vґ�6S�&�_0F�+1d4�q����,�	u�P��}��� ��5-M�6m�7Lk��1%,b�w�'���3���zF�^��L���&V?��ץ�ｦ����=4��m��N���I�����g�������ܐ��UF8z�-���V�E�Xi�	IU[��M��;;�5F��۞��QĶ���ok}��������.�b{�,9����{�v���,�%�Dh�^��ib����CӸ�3������$ciy�6���P*����O��t�[\��������<(���D��m������h�ֹvy ���<�Se�594�4X���C�Dͤ���,�)HT���Iw���}`5Q�?�=B�U	j|�/f���^��q�A�Sl��p7+�_�4;-id٬)G�
"}�A+<{� ~��as^�������8��ͅo��6ܦ�c��G��BW��7�}�J�_J��8o�+ ��,��r0[.P�t��Γ���v�J��(�S��PoZ��"�F�Ϟ��\-�w5��E���F�C�� �':��A������W+&�i����F�bO7L3���*����i��,����>�޽�s��UZ��I�n��[j�ZS�CU�H�	nR�����(X�/��X�k�f!��j��m}R{~�Ph����2�,ږ�!��PvU�*�OG�*Q1l��s�N+�I�������r�$g\h�sYVq�?�@qb�aA�D��ʝcn�|�f�W[�gV$$!]������V�{�Uqw�����]���w�!�c� ����p}�Zlw��锠\� ,hN��4Zt���V�n�'�W�}�	�U�-j����o�t9�1!3X@�
#a��1ٖ�;]�Š�b,�u��z�/�Ď�fA�?~���˽�O_�9f/"�0!zC�C�����j�X�`��O��ڇ��u�,w�]2���j�a�����<:��Yu�ygNa����),���FcxW���{+����jl^�xk�2��ޚ���@�U�umi5
E�gQ>�K���uH4:̯}�-�>�S�m��r���@E���C�zuj�:q�\܉MLA·�9�j��\�=1)���V�
"��<��«K=������L�g#��10��ph9'�.F(�@u4 Fh��Ghhe?Q6��<�����y8�T�5�`�o�|�/Rd�������hz����{������o�+?�a��RBF� �$�k����j%�w�"?�� J4)w���ͥ������g8��l��k�S
'� ��^���W����}O�'��~X7a.5����������脓(��P�Hdhoω�_.�7!0�D�w�jWB��kB���F�ӱ)�����xyq�Ț��<~�Jo��
��	�8G��<�9��oT���7�����:�YC~SD� �����B����m������Lۘ�_�x�@u���Ńm,�˻���!��s��LV����j�c�o��P�cC��`����W�V���n�y�����@��ނ�8%�Q��l�U��j�E�Ǜ�	á�i7�2k//��p������7Y������^��iȲy��Џ��t��:U���}����H(�n=n¿ ���]S�:�%��0>4�/���7i�Wx�TR��뭾�x��K�"���f#
v��_3<Ű������H�!)s���Y\Z���dڀ�|x��y쐼?zz�b�%e[���0�ipg=�����W|�:)魤��M�vl{&5�֡�G�*ax��&�(p�ٓܨ��6��-��/O����N�e��x ���vJ	��{�5���q���"d�æ�mh����k���}�G�������uE5+�Ϯ@N��ЙF�?�8���SA2�X��ɘ6�|�7�Z��!6���g��j~:~f�޸>׵�j�FΏ_�Gӵ�6�r�@<������b��\׾�������R��" P���8<'.���0yC[<��:n�B�/��O�zc�1f;\E�aq�|DrP���j��*DϏ�s��.#L�~DF�;�+]�����j��פd� �3n�ՅøLos?l5�C��5���hnM  ��-�t�oG�x4פ���=^PR=��H�/S�3z�!��*�޴�����;#-�A����^���Ō����\|��¤����`�P��`0�ө�����~�@��3�I#��<�7'��jAɹ��a�d�]z`��� �+a�و���OC�#���vy��fV,w�e�%(i����&*���rz��:C�h'�12r傿�{@�����XJ�~�Vd�h��4#�j��iW�s`VCN[H�K�{<��\��Q��TfV��]�m^��όc��lF�!�9ل NF�5��ԧU��~/Q��������ʱҴ�.��|Rz���5z1�k�����'Y�7o�"�R=�����|_�4��^�+�!i2\��I�����p.9fW�&ط����DOb>��ǓXq�zzH�&��	4x�d������1e�K@M<�E�p�x2utgw�;Ԕ��/�x�5���Cq�{q��`6%^�(�2̜.[���t�ƴ��էO�+��,ر"�b��U����fy������6E�O�����[�9�8����~��}!)��$�M~���hnc�q�v�L4�����p����q�D����Nh�1Ud`ꯧ[py��6Z�� s���m�J������=�����>����6�ΛՃxOˎ�t�+������ҫ�#��ڠ�Ј��w��x<d�DHn��i��g��o+g��m9b���nm���4�����Q,�iba�\�SV	寰��Jb���0���e�zx�+����"8"�M7�5�����s�W6C˽���%P��Ύ��|�9ʸ�����T/����E��=��`�6Ϭ9�
�8 {`��_dAA��Ke���;F��,Ow˅ee�lӯ���I�{v�fFSK+�ʁx�d`�z��}�LM��~�So}���]�l�\�p��C�gW��?�_m�0�}�y舌~�pZ�@������^�^����T�4C�:[P�e�ih��M���݁f�M�ZZ&��X�k]wdQ;����d��4Ѣ��}�͝�ͷF@N���������J�u�l``g҉�ߥ��Pbv������z�� Ը�Y^��Ϋ+��_=���~|{žv�3N�C+�Fڂ�����Q���Ғ��"̎��-n���9�|x���|��H������3x��n�-��*�����T���i���_��D-��w���{5F�=4�4��ض���kT���������Y�6-fU5��9��ן�=o��d�u�4F�!Л~�kH���O����m>�p��-8+��\dl/ʔ�J�~�o/���CԟZm�s�_<�1��0��yZEM^��:�c? �����K�I!�u��#���LRix)��qI��*x��j�T���O^������ȏ���)��u�~u�i����v�d�f[zQ0���q3��v傄"�d��Y��<.���qR�|A[F^7b�?~�D���{�l.7e����t~�?[=�H�O�)�.��,���r?8��^t�p?��;V�{/�4s!`BѰ�j���V"�U��GbQ���k�%o�Y���B�}%a�O7q��Y38�ٗ�qv	\�v������f0�{���ЋY���<�D�b�>GJ�6�������������S<�F*�"��ݝh_�-�x���x����a�5�h��"��`n�Mr�'�MV�c/���^��@��)�6 {Xx��^I�On=6ru���;lY�l}� \�)y����K����<w���)�s�ۘ�-�������}�A�yۢ/���ꂮT�p��x�9�L��@wJ ��d��}�)#n��4�ڃS��=�:�X����r���k����ύ뎁aa�BKo`�~������7d���:eDj=ss�L۲S��BQ��-n�ku㒙��^�s�]�c&�E^W!)S퀽�y�s�5&�'�""w�Ko0��*�$ܑ?���lʴ���mtd���j�Kf��p1���Z}_i�M\Je�w]XX�=�7�J�R��)2I7r��&�;k���H���h�x�'��i~D�[Z�j!����B��F�[� �D�w��e	�'��(�e�jO��6*��+���N��8 Q�&�a��&Ҧ��{ۣ�;��p�u������ԷX�����v������G(�n\�݇��C���k�ϓ��=J�.J�Z��2���d�.bS�b�'����춱��3���k{�v��}ԶY$�$EJc�K7/����N��I�Gu�?���#���R�%
edj�u���㪓��>��ڥmo`���[�ι�B�o����Fq\���T�z�p�t ���Ti�&�7o�u��䄅�9�\[��]���e�ˇ��o��q��nH2�ݎ��܅��f�b��I��C$:�6=!)z�9�s�d��?�܆�W�ܤh%�|����R�Ϳ�.%�R[ØU�����yf�0j������e��j�a�"؋{��}��,膂�` y3���n}m��<����{T�@K�ׯ�5�tb��r��yJ@B^f(1/���B?�Z
�w�V_{r$a׵״ԕ�i�|������a>���Vg�OKN.��G���=%���.>>���J~���ᡴ�Lkk�x0�_AU83�l�O���f���Y]�PXQ��^w~�|@#>^N��#l�����s����3���\L�T+�Hw��z���?���?
�!*���.V����z~d�Sc��9��oOM!�ܬL����vK�P�~Ů�4ZW2�H��jE[ß#虀��ݷ_�T��^H{�l`����k.��_-��"�����|�|y�����<1e�jz`Of�ɮ��,�ͻ	����zv0pߒ6E?��?�P�*���~����~xk����h0�0h ]�s�}��s��ޒ#W�cJ�I���#X��g���R���X�����2Q�
?3�;��pw�#}4&�&3>����sa33���}�"��������Ea2���Uo����l|�Ƃ.��jĊ�@�vG*Ed�os�9�څ�l����d�^p ���g��B���m%o���LZ"�R��u�W~!9�����=����v�Ff�1�So�i7��+�0��6��k����d�W�_*A�i0��O��Nv4羿'm�Ub-\D�Ծ����K�mZy��/ ,�_Td��bj�fxb ��B���^1���Q�h���-XL�%7�)�1��i�������8�l���OOh�\{ ��Sw���ysǀ����Q����gZ^�{��xMT<�<	�-6��'I�;X<��~��\�TY�Mg��Yͨ�J�%�l� �p���$�����)�o������]��D��eK(l���)�&���I���o�L�z}}���	1	��'*�;v��Cܾ��P&�,�9���8�8?}��+U��MF����H��3/�~��f|�&�X�lB@f{�;���;�G�A X��~A����m�).�Źs1:�_c����������ak�ɽ���[�r�\�H�O�}�8�k����ST�a�t�G/]���ĕX�~V�&@g&e��C,�Ȉ�{�Ģ+-Z�|��:W�SW�A?Y�w�J%u����r�G;>��{I�s&8j���jK��&q����ή@��6v�f6f���i|u�mykF�,<(ê�]�4��?�o� ��G�}���gW�Y�I����d.N��:7��:낈�%��`���Q��e%���Tt	.m�z0�Ƃ��ʸ��]旴��G�BJ�I^�����<�޲��mص2-	@?�+��� ���|�{2�|u�>)&
M�`���g�:L}k����-�#�f����k�O�r<�H-��7�Ğ� lU)������TQ
8%�z�x��t�gR���{��}r�4�+KĔ��k�7�$Q�/>�Қ��9W�告����~�UC�	{$��L�%=��ߙ��.��M��Գ���Q����U�@ݙ;:����a���T���B=���n�����.K���[{��nb��Ζ8�� /5�7�8g'��_Zc�L��.#X.6$��XV�Gɽ����?['U�
n:̫.1���q�(q�ynz���Tc�����!���R�ѯ4��	w��:�P�L�:w�(<�U��\!��/�R���P K�G���!an��C�XCJv�I���k���E~e9���B/uǸ��yM?��L�	pq�\Z�aJs�u-C��j�N�1�C��b�M�6K.�Ő�O���Zc�5l�)�T�œ;]��P�D{�y�y5�2w�W�Az��گ��pF/ʜ�X����@����E��u2X~�}ł���h7����IfM��7��<�/G��6$�
E����<y�~��%�׹g�<��/&���#���X�i�!Z�BJ �Ęť��߰�r)�-�뿅t>`Gↁֻ���1^ab�����K�	���|l,���7tŸb�k3؋�F����س4��G���=<�'�OK��ūR��Ox��rP���ǝr�g�{��;<m�k�����ȶg߾"jG29/Қ�I7a�r1b�ݜ����ZN�Ҫ��ޓ��\vm����),��nR�/q@qd��4H�	�f'�z�'F\���TX�q�2oy�����JZA!�
����ի�H���W����/��r�'J+���C��RcH(�u�K[<e!ca��e۞����ãǱFsΗ�-�Ce����q��+��p����5��u��u�8�w��l�����o:d�_�<��y����4�W5p%*3�\�7聍�w/�|�g�άύ��xq}}�����N@'Ͱ- �8zaƓ?�����~Hn,5���!XcY��aW˸H��-���b:15,wŭsE�}|?�),'�*v�w��	K�����Ǖ�l���T$��dq�2�~�VV��ONK_''��uz�X_�*:����a�m!?#�z�q3���5���G��q��k��6�Ć���I1��O��$��G�`Ii�?3P�����_mX��&���F�?�bG{����"u��N��@r��q�!h��������f�r��G,< �=�g��ma�3�a�B�;�J$�z�^������\��=Kr/x���>a ����xo�}��*^��٭'���ڔ(��G2���"����&0}�a�i���x�4�[�3�f���_�7w+�P�>x[S=y�
�7�گ<�!˃�i�n����F��$\0%�&%2����ª܂ZG���g�$��p%��cVI5{ ��+g�1m���#
�O3pYUFXW�Ͼ�=�X��4���{�чxZ�ƒ�hƭzh�I�es�&�l����ݠW���^�N�2J��)Lw�+��K��r������_�]�W�`�;O���-�3U��~4��X��b�M�f���bm��BR�<�[9g�L��r�/˂������MQ���r4�ť����J�}k���o/����õ�vi��?	�� �2C<t��a�j&��~Á��-�d�kݗ!E�<􄆪��d9m������+*�:��V>�����Y�Щ�Tϑ��9hd�7@q-��7Y/��_-�Xr�Z��]:,GFb��b��oS�\r�Vf��v��p�x(��c�r����JC�o��/9Efݻ�������yy��#���7������^o��L�w'�O��"�T���*�G����
�C�'��F��B�b,j�|:�#N]3#�ĵ����=��ψmӯ6��\��X�kt�I�9�~���(5�N7a?{9DuЗ�lX�TY0&��	~��Ux��ֽ7&�0C6�UY��Wܼ��6O[#dd�����	�rZ(_7k�ÝD�;n;���K)��B ��6�[=Eg�h��	��3Ew�o�o�Q$�d�#��v��g���/�����B��̀��z"���d*����5��r�O���Ar��>�h��n�����+znY��[LJ䕺x�*�/��HW�!M+;C��w��y"��@vl9�+�Z�]t���,��:�i�t�T��%hT�ц����<޻t�T0Y
�H�-��\�8�$I/��j�l1K�����'�.�8�8D1>���޳��~>�`hb��;�'�៉w*���Q�30:�#�P���
��p5�Θ�/]0��p�:C`M�����2���v	��ω}����)U��nR�Q�&����T}2Q�ր�X�%�� A����k:O9F�[�d��$�-�u������7x�a�O���l��t���	����E��'��}p>�+�SA�-Q	���:�Q��{���gn[�OD9e�4�@N�-��7����l�r&���݃��q�_�����Nm5���)QzR�z���q��v����%��Ǖkq�Ŗ���u�����Y�Ý���mW;8|�Uk�r?`J/����t�5�!��9�A��=R���jϾ�8�c�ӗ�;s~p:��V�M+;[�����Q�4�5�>�͑�d�ؘ�����BLOW�a�z����r�eѣ�a�����;�B���/�_Ƴ8���|��K�`�a�p+��C5�D�n,9ԋV�����6"E7� �� �|W�e8c��\�F��-�Q��T��&,4ڗ���F�n2׶�w���Dqd��cߺܟ��u�L��90S�w0_׮���e`ް?c>_�2��$��FL�ۺ���I4����a�/���{}UB���$�.\�B�B�vm.4b�nUd7�A�w����In^���p�c�4/#&����LLM�s�*��+m�0VQݡ�b�l�{�y#p�����U&kN���Z.[��+h�&��P�KK �Bհ|��[`�r_�[^>� ��13[\�G�����3�5�qB��������^�x�|���0��z�98�X:�RE�,0b0t�����+;<^ݞ������Q�%mW�A���=�a�+��&ey�T�pL��uj�m�t�]����`F �������ʠ-�_-AE����I���!��ꝫG��k���َ�%p5��9��6��'
��{8��{u�����)�^�TNӰ��Y�݋��:	1�ޚ*9~\��8�8)Ҹԓx*��ah&T20xv��o��l.�ײr�����`od8�����ug~75a5a�~��^5[�#h���Vk�C�p������8M����ұ���`c����z-"��-�)+b��Q��H�	py��A�ok�:6_B�8],>�l�<W���Z�5}��7n�u�(��**�Y�S
�̚��sܗ�G^B�}CVL��&@f:I�Š�#�� �w����Q_��P-�-�D�v>��Bι�h�vx��FZ´v��J���w��9����!q�N1����d�ɖm�6��{l���}������/����^n�Q}�4�����+�M���ye%^|8I��	[��.J˳C5����fdD|Ik���dTdJ�J�E��~c�g�$�rHZ|I=O�@%���ճ��`����d�u={���Õ���k:K���w<7G]��FK�Xx�L�b#w^iLJMH���G,�x�(�/��3���jLC`�Tv�ElAS=K,XA%me�۩w[�ɇ󉊮�/�Y�ŦG��%�yg��@�������vP��ᡗ"�i��Ɩ�f�Y�! �u�Yd;ē� �;�]py��~UN�]�F�n���MM"H$�@�C��|��L��
'�}4��V�������ʯmeQ�7,x$���kYٝ_�J�%,�(yI���|�Da��;�x�G���Y;�$~"�. \��7�#�=��J�'�]㧷���G�ͦ�q7��R�O�n��|j���C�ƣE�dq�\���'�������O.�rum�I���첞��T���"�Ăr��H�$rթ��Y�!����I��V$2
���G��T�YOʸE��w`��h�=X�-��հ��Ų7����ql��0�T(s��q%#���>����[\�M{����>��Q�6��<Ii	p��7&
��[nh\c
[nk�����^!�~��s��J�MN���� �!�&����R���u���	��T�_8=�:^�\����i�a�S�=�MG�N�����ݫ�w����Y�M��<�vO�x���}=�������!�*6*
��g'ڰ�����$�ʶ�sz�}���_��	���(�J�._�ז��~+vCn�z��_�D��Bj�2|+rA]�ƃ�Z�r�N@�>OaG��H����`F�'D�cV��zv\6T��E���t�ms~F�t�=DI9x�ۘ�Y;��1�l�vh���l���D�:�#su�D���,������Z�*�	���X�e�T��l����'����ԑnCp��U�~��WF�_��6ˌ->&�M��/[�,pi*--�U���Ը	L��\lm0=��t(�Դ>L�b�Ӹ��&){�O����6u�>X�SXޔ��������?�S8�tf�S<e��������@�3�ג?)�ѝ��o6	=y����x�'�����ϧk|���'���C"��##;��qSMyyy��1W��6�e�Sl�6�1|׬c.*���:����-�D,�t��> .�����S���'��5̜]���d��x���c�u5���+��Ë��EI��~n&k�X�k/~��Q9�6�3�F���M��T{���ԤGC�]�^Z�r�;~�Rܣ�ǐ���_7�aċ�X�j��S7na�Mvwy�w|�s�>�[�����Ebff�����őL�&)�շ5� ��f�<h	��,&`��Y9��=���x~y��-�y��^F�y!J�:���>(7<r*���H��������d0% ��,�pC���P�F/�f��+��a��z_��&pP��U�qY�I�/��������J����c4�93a~�}�Ō;8���;�p�/z�M�&�uч^�������>����{AsːG)�y��۷m��x*�**.{bZ::�#0����q�rL�] _^�_�6�_��ډ���T����ߊ��qb&��g��W��F2��k�#R�h����?��8�E��y�i^�L6�BlA�y�<�}�K�[�Z�ƨ2�'�pE�Y�^탆�	��y��J�?m��ף�OXG��^�F�6C��ֳzEEA!a ��>�J����9��i��PkO�AрU�UT���(#.#�Zw˙��%G4R��y#G01�"n�b�?h3�Jɰ�v;�ִ��=֍�.3�G������i=�x݋v�=>��ݶRv&�2`��g�}⫧]����F�8�J�u;J��$�.��2=-2)�g9V֩u�3����GI����L�o�\�8�u�I��.����\��m��M���g~w��d�E%d��dڀ)�M%����t> �S�l�������@,#
NdŸ���v<�d*�qQ��M#���-k��Wd\��O&�/���<.Z"RW�����F��� �W][��Wx���e$H'�T
�s����#�v%c�pct���=|��`�����Wƃ}'�y>t����,���n��b�o�ESc�d�|�M�z&�oii�Kw�=a%9�Û"~{(����K���(ْ��]{a�G^�ˌ��ͅGhC-��@��ˌ}Ï�`^��^���H�N�O�>���9�l�qC!��~'����"��;:Q�zW�r�ܼ�#�����E����K#b�`D�'Q�����Vx��Шk�Q�N�������H�;�r��4|�a�#pB�xE+�����o�*�<���_���⋷^�������XT�/�;{���R0��D����\�k�T�E,����s���:�L��YƯv���m�8������ѧ(���$+% ��;�CڹSr?��mo�G􄰲�6?�߭Ơʾea�'|���>��[�q#o�+���no�)R��O�~,� 7�A}���ea������o9���3����MO�����bPt��B����}�3�؉Ա��5ރ�9�$���u�CZ֒���e��q�t�=z���}�UQ��/�8j��G�|^�C������7�^d����I��JN7_P! RT���$����$�L��Ҹo��\)K�������6R�y9yK���֗��4�Y�3Q	ɹy�kV�T�eX�[�?L#!��(��t#��ݍt��t#  -�1RCH���R��!�0�������</x�u1{�����Z�0z����D�	0g��S��xTN/��sO���_���%��_mcJԑ���X�N�a��ٲ��HhX2��I��@�) �)}[�AFۭ��kvf.!���Cf��ٮ\��t���ɗޚ gL��&u��Z�q��,\�����mi�B�>��Ij�H-�(�<�rF�Z��aj[�Tڗ�D�S��;�F<F��I���Gp6a�A)NO~oV�����Z�t��Ѳ��>�vP���;!��)}���Ǡ�A��D�cǏ�;��0���%����WrC�����$��X�xM#P���ޑ��m��0�+Y��g�`M�}���-6���H�B��}A���.�)�.�1µ���$�>Z����%e���%���BA�丂^�T����
"�yo��YܢN�<���rÔ&�O��s��{�fS�}F8� �$-&ZD(���M��蝄j+%�w��N�#���I�l���0>���Z��=�(�_s��~ �d��2�C#��sh��?�T+b��_q���Bl�r�I))6�}7�K&��=AZ:	S|�!�6�" ؝lO����V���Nm*�F��P"�����D�xla�naI���Z_2��D��CJf�}�6�/M2={��h+���P��wgdA�jY��{tV������S�\_�ם$�[_Κ�]LⲆ�����ҫ{����Aǫ���Vm�R�{�%
�n��w�w4�������b��wM�L�h�8�g��"M�8�ӠT�	�*�v߹�UZ�<Cn�uy��wa��B�{���Il��т�q���6��Zoy~)������/:ӊ ��w��X���dX(�}�w>?
�Γ xq�����uH*�P$6�B��tR׹�v�*S_�����I�D�>�����R���3��r%�6Ɲ�@�KS���"������ə���-�k�P#<<>p���ycEVX�#>��pk2ʤ��L~�Qo4^�v��� �����ʬbt���²�`)��N�Cx�kvO�lcy��@�k0	�C��Vt�H=v\���CK=�0v�jJ0���k��+��	ӂ��2ؘ�~�D!�n4#��6��;&!\vĈd�!gp��#V(�h�5��0���Hz��'B3�+r�F_��>9������� ��-Δ�W�����ǅ	��N���������	�p�f[��&�T�;�_~�x��;���3j'�������Lac�U�ͼ�}N �+mϏu͖��A����Rm3�B܄*�Ǎe¹�e�o717?�>�_����c����C
@V�K��|D#S�̌��J���3��`��._�W폞-����nX��D���'���\�n��bͻ�?��5�?�[.*h�t��֖-odK�)�%-�:lJ�6��Ĵ���4�g�薪L�I<��}�B�A��s^�Zk�zE�C���0��/~�p�z�V�*��n�S��¬�J�Q�����Ќ��!�p����ö���5�4�%5~F�.ܧ��ݏ���ܰ/�+����ݜuRSU3hi��B�v���ym!~��Cu�X6���'n����6iPϽg,|�E+�WZy9C��f�<��x�0nQģ[;__��Kf�������&��Ć88��&��`�D�6����5�ܰ���Ү�������h�p+������1`��[ʡ��MwY�SK8�G�xKZ��J���	Ji��oC��Xp܀ ���#�2^�t��V��[3Z|m��NҠ�d�(T �z�;���;d����h����שWֵ	0:U�5��o�����KzLo[N/�5F�`棵����E���Gy��y���E�'&����0/�U�_�	���޿�:T���,a�L┽:-Ҷ�HIK#u�hE��8>Ͻ�@_� ��GT}P@ �2{**��b��'����/����&#�a��6�ؓ�:��tP�ն���U_�x�6N?f%���hXz�bL�\ŷk��bǁ���T�˷��f��������ߛ5�����pt�$�_J;l'_��%E⓾l|w�x�&z}+�;4�s�\ƿ��=ƛ_myR��P����T��?ko9�~
�ǎ�b{S���FE�Ђ�f�JKK�W���`���}]g(��'����A&�{��י�i؀��d����:�1��:V�2��S�Db�d�	��v�[(yg��J
�t-���'���wD���Z2��|":��>�����Qg��6*d[�'�Hg��PS��O�^Ćap��� Y��b�^K�䷟d�Eք������VA��e��G}��O%%��4y����?$�g5��Veى����gi���t>Q�cTQU;�Hb�� ��-'㐤���|*$B�/��<��e���d$RL!E�I=���pe6�wR@ޑ��a�p���[��
}�$��o����5k��@���_��Q�p���0{�*�Q"aH-{-�T�K�=K�#�����%z^uj}��u�����ЖE,���3dqc/)�^�Q�7�;��߉���������.���N:��^�f�G BO;X����]��./�v�h��soP����'�;��lo�d��:��$	qh�y��L�	����?H�o�ۑ6��x��Rc��ǃ���G>=gq	-��{��A����ނ�[jē� �T�ӣ6�����q�J�FX��ף��fU:���?��w�sr$��]��d�B���J9R�?�x�k����`+�������ǌW��`�j�Q��a�Ɣ�Y���[��8J�O�� ކ]��ԢR���7E����~2+�������I�Nr��O~u���O��ێS��IQ�[�E!fs��<�㎊���H3){��&�����L���x��܉��>�	$}�����O�1D�ͨ�IU���zW��{�����2u��]O3��u.I.Þ��+�KPH^͸�q������8�Je�9e�d�����j�[��Z]�ͯzS^��g�F-:���U�X�a����Sfp����
=AYٔ	7COp��W�d,JJ���r�T��8����:�WFc\���sr��oz�MY;?��L���{��u�7��+��L�3�C��G�<����寒򵎣�� ���w�Y������w{�)�GK���R�D� 8_`�c��Q�o[��r)8��M@�3�������»���� t� 7���1�������fB���Q�����@x�0�߳��|.�,hL�`���ME�B�	P��{w���V�j�t�X�j�c6�[�?|��֍\�H9�Vs=�	�	���BM/���큖�;h?`81VaTZW��M����T��.�ݒD(��0�盰�N���X�>R�Ѱ��-�6U3�b�@�*R=e�<���~]���05��wFvw\k��2�5k��V�L$��~@7����j�]�y������Y��������"�66X�&���MV+�u�L�2��k�Q��"�6vv�����@(�e?Q	��񉐭��J���fS2$�eÝU����p�����q��k0���	ц]�����<1E��{n�	��Z��AP�s{� �L=�b���rW�<��~����>/�u�3о;9���3.�:^�d�$��+�9��!*��4�Iԫa#�k<����7��j0��R�:C����7�}�X�FF�$���f���.a0?�Z�W��
Y&��3/���jQ�KR��'�Mq�~1�}Y�`'�OX��Py`������2��/EC���W#������@VG�5y{�j��[<��}4yQ,+�_��L�;˦*���{(7e�hODc�R	���P"�O�!�|+`�7h��o�w�!=���.s�4vǄ�!ò��(��OL��2Ѯ{.a���R}���fy;2ݴ��e��[��l_��b ������D)/�e6�e��zT���آe%���q@Q���I�f�WQ��?ߵǔ���r���$%���9�k��V�d�w !߻�)@�����~���U����m���o���fgz��7��3��Z���"qta�RR��I###t�H����~U����'!)����������{�)>&�᝹:c�FN|2y�3p�z06	����"����B1̒y|��*�H�}���o�X�d���6��Ï˥��Wo�zuT{we���<����d��gJ:Q��'�/�"^�kf�N�v�c�+~���|*����^<l����v���.���m����dz1��Oѳ�'���]V�,�\���U��J��$�W3��5��3E��dOP���x�sV)�Ϥ$0;�yn�(C!�Yp�WN�t��=
*8|u�<픤o� �y�:��Ȩwa_�!^,�׉kp� ������ry�8��%�5�
���\:t�����R)Ļ�~�&�bT�L�V�"��_^h]d袞�Iv�S��B��Z_�2��#�>א01�mX�k���g�=+�<�p,��E;��@��w�����¸�/����I�O����k:�H�!�xZɀ��|�@�\SQ �lmm%db-�������|��\X ���f[�Fyr������#��V?�Lv�@o��������݆��a�{JL�tFz� ��Lg[�'����NN���M/��k��2�b�7t�h����,�E��S6��Z]����<klP�>v{�8`��=��O�E}rp�n�_�S��{�j����J�/B�iUu5؇��p$@�m-���I�)+v�=�X��Z�'�0O2s8���D�K���ۓ�m$�*�����F��O_z�O��\�Q��DI �* "�4H ��qɳy?^���]!C����py�uǽ���%߰^!QɄ��[[�)��ɓ�I�����Z����~5��4G�j3,��t�t�Y��O�F+������㟭k��cSS����a�p[q?��D3����+��Zfe�+�Z�fD�w6�s�`�a�[z<#�:�����
o��G�_�����G��#�Q�a�m�b'����%#�F�1�]*�)����A��'�!����0�����`۹)�����������7�!����]���*\h�U�)A�ɻ/e����l/�׫�����@<?#EUE�9�jaar�yy2�� --X�P�Z__���.�.��Kk����{�臾��x(|A��6�B���e��{���Ĥ���-!���G&��m/�_E���u��;�c`q�LM=�j��	�L����� K�/�n����S�s�ڔ����O��7�*$�j�!d��	�w���aL��'��,����C���O��c	5eN�R��D+��-�3%u��WM�\�8�F:�)z�zwjy1<����U)�U��9�o�����~a�{���y#��y�=�~�'����s��w��d�2V�9Lw���^Q $L-T����]���L�j�vޭ9)��^�P�Y;R^=
���:l���z������I��ex^75���~�Jb���������<0�E��O��{��꥚���ib\������;*�g,��\���ed +X����.�5�r�W������G�6��������/�R�G��~ɮ_�sx����0���d��r�@�6g���0b�h9����c`*�],��0�����3t]��#{w�'Gb����;��-k[eb#�4����\�A���gE�x��%�j��N\�������RM!f��&@��7�<�$pK��b��-�@xM�`V�0���r���崸�R�SO�1���y+o{��)K�����O�%�Nm�+E�3\dW�kΖ�i�=���=�n
��9d��R�i�jJ�r��Na�4��U���"4�#DN��9�#�krr=Fee�#�9NAA�Q��`Gb��L��ш4;<$d��#@�	���b	�}�����e���1�g2�)T�L��HRRk;'��r�Zh�0��<<2���9﫩����㽰;\ � pѦzu7��{m8����w�I0��_Ow6�=ǎ�/�l��F��F2M��p��^�ojf�^����mc�� 	���ڈ��F ��Xr����!��Px�/^�m�;�r�ca ^�� �<a�,���f�m��+ٴ��b�yMW>�xM{��N��HĐ$Y�O+��ɜ5��T���	�.~��S<t�%퍤���}����6_xmooW��3�AX�Ɔ��V�i>[y����v��7<|<Ai����7�4�h���Oϲp��jK��@��u���!;+�/f�/9������=��oE���>��ND!66�c�`pYX�-����.©�T��[@G\�d��S:F���}]����U�%2�5��W�:�`+�w/[ـ_�
'��G2�I�����͕�V�F�%b�Svo�agD$!a�0l����ޗ�L�z�$
��<\�{���!mԩ�F�93��|����T8�V{��C�]/��?۰�T���Q��B�LYYa��+�B�jy����T����M�G�	�#��֝��Zm��p�9�#�>G�wn��a,r�bs�X!#�=>�)�m@��c����%��B�����a� ���>�����)7��3���n�潕�k<�6���]+ߦ��O�Z��55�8�)Ē�l2��P��m7mG7��Z�Q�ЅfGRIIɲ��ψ�'E\D;�,b7��F���u��5fTy�^ASJ[
���]cϢą����5�9 �׭[�ݲE�g�)>dgZO��V�s=s~��_L�T�����w�K��R1=^DMB�1` ա��:SZ���S%%�|ji�z'�ak�U��}}F��el��;�"�D�/SI�~�-�������,���KD�j�}���
�ʕ��5�x���qy�O&�	k �v���g#��ԯvK�0O߻g���x��(Tl�U.O��W��c<{�����ASzG;Q�8�Jdo�}}�=���3��W����>��� T7���f�&`Q�/�]��"���8T�* {�E���Gc�f�z�CO/�>xv��/��8�{�ZUt�Ҍ&{:4:�ibb�>�TY����|Y���6*���-O�p�wm+;;��EC.�����45[UU�< ��yx��%��Dd�\��" l��E˙oqs3��R�M�K�E��pB��qo����s<tr6gz*���=�{����Nm.��W�L
#�Ap�D�1��&�H������㚏�1�gQ�p���Y���W����ܾ�Tl<C5�}�
�ׯ�(ʍ��C}�GU�|v���ztG�]f���i\O0�"���6�`�KLW�Qn�βC�綌sn��M!O,\�JDWk��R�S&��-�7��>hu�=�[�Y��&�ޯt�ȷ��ҺNgf���X1�s[J=[j5/̆� a�0���� ;�Y<X��8��ώ����T��B�;+T�[�`�-â�&6Z�"gqf�>������a�������Y�p��� R"ù+5c����c8�&A.�C8��Y�_��+�<�M�!�����@�p?�d)��.��v���������"N����j"�]�⌊���;;���I��|��ݩ������h���SWG����5`��Ğ:/|���	�;�k��#�3�(_@��B�@�u�����Lx��nq,y?��ο=(��6��iJ4�0�dp�.��Gk��\Ȇ����,ߣ���ӗ�o�L�n�Ok_�/[��4$ y�0�NǃZ�xR�������ӊ�f�.'!�{V������Kl������W�+�3��T�;/�魥X(�s7�yl����������ؖ�ص���,���n�w~2��U�����cXHt���
���Bd]uף� ���p�h�D�_B�V��m3[����OԎ�Q��������X��{�7�r�����i$����=Q������D�Ǜ�+D�f���;�lV�L�
m�D:xV'2�V�W���WC�����{�w���eb�/�������,y�0O��1h�Dʟy�(o��C��M���S����p�0��nQU�!pR�3f�8$?S �Y���_+�nIlf�o��B�"|5c(���_'o�aJ嶚8�N�9ԏ:@>2���(�鷰�8�z�����[m�7}�cr%=��k����Ӣk|II)F]�!d,���w�+�at�M�s�.2��5���VN` <t�pi��soមk[0����߫���ҧ�_�/1Z�����K
�X�����!�@~zs;Y�]Jŝ�#G��������i��C ��TTT����WR�'
���D����k+|&��L��f���M�ϵ�8�ͯ�04�Z�����l�m�x�M�l�/��^fe������;�e�\ާ�;}���z���i��zB���?�O��z O��Wi!�i�}V�c�8V]九-�1�_'i�Lj}CA��!�;� �}]%ů�\�Y�=3��9��n�j����Q]�*�����G�}�F9C��q }���T.AF�'ȃyڃ�p�_�F'���O׮���Y�r-�vҠ|�3z��&,%������J[3�IVN�8��b�ޱHh}��n��dG�u�7�+}h'`&��հ���SA��c�R#������Z�@\�&�g��F�c�[;lv�Uƾ�_ 4(�B�oY&����F�:��ޖ6�ܖ7E�܇:�M=9�ȏ���`�GL���T�9tI)��M.����w&���F���nM�u����x���gAPWbA�e�3_�d[�t\��O�c0�y��ɬ��T���g�j�M���Z�P�������Y������X�`kW����Ŵ=��v�^�9�z���u�l�R�^ژ�����%�U҈��d�#�q���n,��oP��G��ƍ�����j���Eg�n�<aŕ� y����c� `���v,���2����&���{.K�E��q��'F���2��8L> �p'*8LqN���1�*5g_Î���<��}[���
����,��=x��1P�&eb���[y������`{H���ac#L7����'��饈>����.�XTi���Sצg96yz�ƓP���[Խ�>o֯{�`pi_�#
��j�����\ScRXt��6�s�=���$۾�f�8j��SƸľe3�F��Η�S�Ь���"q%�?�@yE��b�B5 4O���IBϥ�Y��刯`����{���U���� �F���t���/l�J�قf�^��s��2�L]��H����/o�t��|-���(L������дq�^��4�U�?J�gy*�μ�}`�W�|5zKmcbc�Ng�ĩ��) {���p�r�i^��:�=��9� ��IJ�ZQ=lԩ�<��>�pʯ1'�b���x1TSF�O�3��)��}�kОM�����R�?��'/t�r��7Ęo���S\�ש ��E{�ԯ~
{�����w�@���G�2��N8X�:X�"���'6vKO~���U�۝�d�^�����)�.�d4�o��/��ܖ��'�^0bE��e�[��fl�!H���7�ӏ�[���z:n5��7M��H�r�vk��;�����{��� 'Veoo�����a�_O%&|�9- ({�;��^�v<*��{�Z�
S=����ݓ)���n,������Y�ۻO|"���AE�WB!ɇ�h��#��w���c�ںl_Ӻ�m�R׶��@?�ig��%G�X��U�pG����ZK���#+?~Q��S.� ���AS q9.dH�����H���ݛ�o���|���@p�,I�{)O�?DN���8�I�ox_8�0�=w7G�eevoM���wM�x7>�W�<�=�Y�������b��'�grl�,2(�3��::����c"��:<�yF�C���o�0]�!ߟ�\��	=���!6G�/�rFq��Oh�Z���a��TG��g9sT���[��9��Ɍ��*�rm�tC&��z�[���a`����	�q�Q�P��)���|�k��{�p�6�tg�z�����+�`>pw}�
�z��gNO�z-A����>��HtTvR-�n�� �j���Ĥ���:���m�ٖH�~��8(���'Se
R��Fz�e(-ZR[$�YP��`T�I%�u3P>Uu�2,��xb�_P$��\���U�A�N}����&�/�>�a�Y	:*��Yy����kۛG���(�¼������۷��JY]�l�9��h�|f��&��Y6�2�wq�8���ĚK�"\&���ߩ�^�������=*�u��N�E]�E�@�����ͽ%>'�FVo|�U�{��o/m<ݲ�_�Ϩl@|�2#��yĊ�v�N��!���:���O�Nt�4���Z�\����wkFB�Н���=�;�t�C���E�C�����������:mtz�Ɖ{���mh'���C�\7��Aq��wؐ�������;5���y�\D�?G�kQ!�޻Ab�6���j, t4U5	�(h���_���	�pHߺ�1����	��Խj�b8r����+z2�GEA�p�H����s�Xs]��}�gR�mPG��m��s�n�B�������ϟ�m���9�op��$.�y����ָ坠L4�Fx�e9X�F�hq�ӈ��vɴL7%�v�/Ci�� �~>�-:t�^d�Q�HS��[ʑݧ������_��B�8��i����Ȍp�黿��^`���N�4�VR��U�#ď���8<�)+�vIe�O}=�q��8,���A��#�#��V`וM�xH+#����A�R��z����y��L�Ċ��]4x�9��ږ���uG�E�ތVg�7��8���$ r�螯?{'��6�|;[�cP.��(��h��/�j�oku��
d�T�}����m�����3���I/M�{Tz��)�?� ��3�Q�-�Ɵ�A2���i�
� z��)����PMOg��&I�a[/��_��g�|[,������p�.6!�Ch���x ���D�`����B��cߧ��'s!O�{[kʩ�:ɞ�=/	\���vJ�����M��}b����z���ug@?�NB�ރi!�ߖ�U���<g���v:���/�m�݌I&�u��充[|��0)�4��(�~LП%Ŏ5��F&?DxG
Lo������].{p���V���WٟxcX�j�ƝTQ��b� �П�X3%�V �3�8�&<Zk�D�,���l�uT�{rd�DY�� {V������2���|N]�k8�u�(*��[#�����zqj�&��a2�y����isr��W���Ϗ)P�1e�U�����g/w�?����LR��(���2d�����C��_2�Q��T0J	w�h¼������~�x�v=24�r��EC{�����w.��{�P��������+�$���Y���ӎgY�:>��ue��¶1՛1�"�^���%\~Ad"�7]#�ȭ(���	1��~ݴ;�
�ZI����5��]E� ��]'6_X�AY�=�|U0��d��:���݀��i5O2��O���[NE�ZY*8׎��/�:��a�
����WЀ������[�z�O�SLI�w�}B����c44vx닐r2/�Z	5�*�^R)~����~�����R�=�G)q���o����{���=*$��_5i"�7�-%goܗ����lr�KN�����Z ȗ����t6M&���) Dǰ�U8ER�-�`�ߠ��񫷟o�m�g�Q�2ӳ���8C@�AA�@
z��H(s�Q�W0Ц��	He�� ű��BU$�Z֚��U@���_<���p{�(���N�ޅ�CKwO3�G*�1W5���A�&E�������)�������kL>�D�,5&��z�{�-6�^�>YC2�w���,�×[eP�mfoǢ�
1Bd��:��?���~L�OKVnؤ�U�E]���܃m+s�0��L�<�����3&�7�i������Ͼ�x^����j�&k]���|��>$h�+y~мS�qp*����T�@�m0:JЇ��2���[��)�kM~���B���yG�M���M#�����B���(٭-�ɋb�e-U?�{%���V��\�.=;��m�����2~�T��~<��L$�g\8���Z^�69L�M��c�B�I�]#��!m#�σ��)3_����vE�lk����q8س��jV{�\ʱ2��+��x�.��������K{�Iar�ĝA��B��1���l�_H�+�ф�곲^=1b�`�c��_������6� ��/X>�V��Uv��-o�x"4����4���&)3n��(d��B�z5�>s�za-�n���&gq?<�yI ���ɳ�#W�H}v��p�V��i�W�_}���99��n������tϭ�I�{�~��t%+{P�u�V/M�t��4��w�������S�ᢹ��b�4,�S��^����n7�鵫�R!��?��M�|���Jm�Rf06���{C�s�4iD��=d�6�|�sص�T|f�Yh�ޒf��K�+ف��|�{�O5ܡ"�?uv.�߼>h7��p�Jr8�Q���<��$����i�7���_��J�E�ռ��c<�	Y��V�H?6��5� 4|�$s��X� U��#W
�)c_t��8I"vū� ��G�XM�쇮Qoh��\k	���;��Q�.���@��.d�2�߯l3���e�����UkM3*F˸����`��wΥ]@����G��;����o�Lw�������v�k�I!�1���;ˊ\�hS��j��<,�R�p�N�e��Ƈ��˖R�0��!��}��Q$��[���Z�y��ҭ�8�r}����0��mʤ�@y�Q�/Q� ���q��c;�)�9>b�gP����މq��
C�l~��d���d�i�6��W�=����m��c���Ο>|f��ܬ����_���7��kDav�)ᵅ���g��BBdzN���h�ke#�7����m�\c����F)��g��WU�(�'��:��+;@4��QK>�[^�d�Ur'�l,�N���mp9iߗ�c!�^lc���E:��D0u��@<eS!j�o�0L� h̀c��_91���	w\��  ��Y�H��z='�ZH��n��|Oh�`nr�yr��^�nHҐ����W��*^A`O�l�Ƕ,�pCyEMQ ���~��5�կ~�Q\��[� <!^��a�y��|y��)�b.�.-��"?���%�e���z��� 5���V;{~*8���
FBW[��S=@�3J'���U�	��}��YZ����0w��l$t�y�q�b�>�B�@��X��+�m��}]T��M)X��K���r���h��|���Q���{��g<�ʝ
�k��A�>7��)QN�V&�ט��>�N���C%%�)sn��wk+|чK|�jٔ��f.�J[�ЎUe0��a�������>n�q"���pws�Py;vwE;<2�-��ϟ�^_�ȩv�F���e�O,�~�������#�ͲX(4*����k�"�@���������f7Ə�K %�G��jumF�/���3��/;s�Hŝ:N����|,�/��E�s���~�?�����ō���L�4l4���L�Vq��t%��P�q��W:`�x[q��.�&~dY��yՔϚ/IL��5��T�x �"}��/^�����.y�%�fZ�s\�Hp %�	�>,��Z�yk���ׅ��2�4ǡ�|�?"({>  +a�=q��H������P��zJCf"�nj[�5;�;?�J(�m��ƫS������?1�#�
�#����`��+��G~��5|!2����x�r��Tɱ��tƍ
\8���lw��R�͢���є���m��DVN
G�;�kg��q�	�s��\/E'�(�q�RΦ=��7Mr~]+G���?J[T%�7n��{��$�3e͐>�k�q����7��b�2����iW�]�(�⠳\�m" ɗ����߹�7Z���F� �+j�(l��c��j��L0Nxt�4�`��o4q�ڦ>�¬�q)l@D@�FqM�zA֚���(�\��eG:�{վ��30��Tx�{_p���wE���X�*(q�kW󽅳cU�r���ٿ�
Mʞ��*��	NF��`������F������dd���n����eP����w�S��߁@GQ��:UW�����������)	�Z���x5%bfG4�5A�!8CeN�~��?�z���υ궊2P��;F՛�7��vN�����<�����L��I[^q��tKATv{���'[�iF�i�,YF���`Sח�ɏv&���rOt�X?��aLa�t]*d�l0Zv�W��A�A�L�L�`��:ڤ(P��~nE�v��1;�&6���J��r"
�`n�T.�u�}�k&Ch>�*�k��e�U;+EqS�Ǐ".B��2?d !BN?�;V����2y���W���U��>���q6�qy�1���<�\�0�n�aLaWgv�q����9�����.}]!����\}r��)ͣ���=��j����R��	�V(=f<�k�fA�n��Ι.�U�D]^C$)$��o��{_MlL�dwJ8h���F�jia�mu�j���Z�2��>����F��^`�9rPӇ]����*�
�1]B�a�������Lj��f�:AI��ON$��6}m�&d��
�u�*s������cb� Qo�t�����R��$�f(��Aa���o�j�+M5�*�oh�U�g6��jk��qZM�?�f�O���M�������'�F�s�Y7͵�8�_����jܶ�V�G���ݡQ@����������h�6���>���6�={�u}2�2�K�U&�����bE��F2�%�.�-W�I�Y��dDK[�֭��1u��r�u��Q��և�||:c��/py䵚�ij��=���+�A���]'	��2��#�krX������e�_���-����u�,!m���(���(�����!R�aYki�kly�'ü}bT�������c��7u�'��D��	�ix%��+�Sk��&� )�f�&�*(&%�F?k^�HD&�Y3B�qtys �e1���|n����®�����o�1��+��;ٗjj�{X�c�⟏0\���)^�T�̗/� ����rW����Q�D�$�n����}���m����D֋��O���k������X6�����(g���<�����l�]?���4��O�X�k˶
��0����E��q������?Ǫ��C^L�엔����FU-H���y��thp�?9�W���.��B�>o�qb��������j@�f�p�]A�� DC�����`���x���ync�z6������y�4��_.ڔ���{6��a�8"Q�L��#��/#��Q�I`
��g/��������<q�I������������^�a7~f/�g<�Pƽh�=��-������T/&����u��z}�C��J��'��?�+���#��o�JT>e������m�R�r�[�}U]MU�i7���U떕d�&S�����C|���~�T�]Џ�?	���)�r�7�4x1��������~QD�yB��i3+�fd)��C�;�	�݀E��,i` �s���{i��7��?[je$<S���cY�`U�׿��*׿��c��9��*{�aV�.!0J�g#�L�V��c:�G�**\��(^o��(�հ�US�J��I� uoE>�	�F� ��f����ui�h���o�q"ZחE�h��ZK�΢+��&�������T�-⫔�1k�K��S������>��78�lvll��'�ITܔ�u���}���TK�fvl�HE@Q5��d	5
o�d����5�kQ�֔�Rq&`)��mT������ݗ��u��w�{��J�q�7R��A����X�7%�� Zz�������2��8o�ɻ�]C}j Ǌߋa�hqF%$$Ե�+<
����i_�wIGU�\�!^ғ�M�
{�~0��uB��඗+����T��a����$L/g�3�a��X��� FھokZ�N�n�K�A���$J�v\�n�l�� ��KGf����{��2=�S6t4���u��Ń6>܈2��t���~�<IBdtt��،ŏ%;$|����a��'#{k�@JW�C���غ��?  � �a�Aʹ�R�1YEPX �����K�6|��A�f�\�G��J�����:<�.@��-^KpY�%oou�]ng�&�����w'v�ݿ�'�U�ї�CA��?�[�/%��.�f��^amc߯�oŋ�ABT����15%_>2	�3��`�h\x������/��;^͓������ZJ=#��\��8NK��`oio�h�F��y�+�8Ō2{��"5Z_�(%������}�d�;H �ʞQj�M�;�4���n�Q_����a7��~��|�3��Ia���\���ݻ��Y~�^��✻��W�UWa�ə#�\�ee {zz�V�n�>����G�)����i6P��	@���T~m�BP���ؾ�u���2+`#n Aw{��;���ш_�$2�W��+��X��!毷V/��uK�*q��jެ��費-���.5Yc�0JF��-{1B�
��=|EIIY�o������@�:Y�U�<�Ƣ�m0�2����CL�Cp�mlR����>௦!<�����y�=+Ǵ�QE���zd�� c���:�=��9_�������G*�H}���q��������L]��͹���l�|���z�k��~\���¯�uݒ>׏�;��S������M��ׅۢj�ޔZ5kojU�Q#j����U�gѢZ��,�v��{� �.�D����}�?�~����9��s�9J=_
��q^q!Gf���*Z�_~��W)�CѺ_�-�&$$+�ᨊ�<��i.��8Ǵ�����xs����E{���G�Ը�{,�Խ6y�T�D�W7d圣KA�/���[Q�@��P!��b�Dv�|��~Eyu5"����ۯP��ײ��~����K���Ŵ����觸$6��½(�5��pu-Wп;0<� ap����ϧ��e�Lbu�v���ͺ���e���v���X�#pBh�zlNWق,����O�|�G8
�G�9����Rc7����X�4���uz��Qg��8L�:��*��N����p��PG껕�3Û?ĎX�i��f�"K?���m�J��cLzx}�t��G���2�q��L�-��7�_�PG�����x���0�~-,Th������\���SSs�{'`w����b��aT��b>J*����0g̕�>�es�zaR��#�t'a3�j��N$i���T�mG��>�l�yZ.�� $��z�*�����s�2A�#˕){�X��9]��͘��d�[OHO������AU\�ԁ�I�e�v�<$����2?�����9G�A���R�:��+-$�^�X��������7t��N�v�./���!gڰG_>��>RF\�}�.Q�u��Ӣ�><�&�����a4��f�����KV�l}�TCBҶ"�la�.(�nڤ��%+�n,�~{
[�=^7a)D��L���%?���;}�s���yHQ{E�D"7.��lc�T劌����=4�E4����ަ��>m�F $�n-P� ��c��!�b���r�������)�g��d��~�������踮gl�Z�"h�iQ'R�Iԭ�Z�
H
�g�	��ҥ������7���_�/E��͊��\Fl1%�O�Uf���gS6I��[CZ��}je9.�S�����J-�P��ƛ.�(:L;��E��J:����*�X��^��x�5���Zb�e`U2�l)���T�봸����c����O���/`�:�z�I��������c=B橨����(����g�Wxڟ�$�/H�gK���ݘ�Urjm�L���#gu
��m_��[?��|��[!hZ=NNi1zq��|X72����"y�*���K|��@\�t��?T1��	�s0ӝ���3��'f/2�}g�ZI��K�2�/C�V�"r���d���#l�d����P홍��Y��lgL	���ψI1t^��z]�^zeQ��,!�j����(�k�a�,V|��˨����Q]
� �N��C���*����S�D�����	���s�Z��}��ɟD)jG������S�&�}qs����y��3�
�.���'�A4h����`�j[�k����±`�E��M$�d.�R�����x��B랉S��Fe|+z�����lڂ:E�`�X �qa��g�&�/;���~"/Y����P��{�w�8��fk��yB^N�z����������u��Ie����^���D�����?��66��L�sb꭭n�c�ЪZ�oEd#8+��oڭ��;(��&H̀�;��O�T��
`Ig�2�#J����H��Z� ܰ��:��%������[��z��L|�#��ϫ�N���%D��{�y��jIF����1����oEzb#�l��:�6q���>\�_��`���ߋLD���nC��uk��0�O��.J|�U)J;#n��:��8Զs
���r'ӑ'�/{To�iڐ|���������!���xGT�秠��)~o�DV[���}W��߈�k���1�����sttD1���E^��3��X��y��X�=Lc{�K	��Cvs����#�輻�3;���j2�>k�����`|h���Y2s����KT��+��ȂuJ�4-�[��$Ҍ\j�r��O]�]d�w���!�XVyZlEf���'\��L=��;�q���.cOg���������Oš���.�-��̜-`�"�b�8b�C���q���C�4�B���8;Z���;��f�烼WG)�+�ߋ��L�o�� �<h�{�Iԅ
����cS'w°t�:�N�tu�@j����xsj^<R����D?��� ���W��Y�c����o�'u��
b:ְ���C����۫ߥ�)̷Ǳ)���ψ<�޼���WYƔG��C|��:/�|���U1��[�������8G�z�����o���F���C �J܍�]�
r����F�����k�>��
���'�*��-�J���\&���<��OM?,�38u�e��]E�z�o<j���q�<cˤ��<{Y�]��y���������
l�<���#z�̼b�.�*�x�p�����,�|rK:���:r��]2�+ɓ���K�|@@������S��X���co��j�9�.s��r�)�-�ފ�12������6�a�>������ǫ�v����^֓���K5KtV�������}�pY��?��	���_��y �w�ܤ��.4��{�Zyؔ��ύ0�+��	�<���jĥ42�X����8e�$��ڕ�n�?�l�-%[���֗��I���g.aN�C�_Z��J�Ը;�b1�x<�O�j�e������(�]~ki���WQRz��[�)`��q$S)k)d��|���!gD�0o<]�dwߒ����f���&иf�ēBpڂ�{d���o��U������"���=@�}	��T���=
�s�a0.�)���Ϭ�E(�CNc	�2�ٵ�}���?���:t�DəC����nm�K�<F���0�Y�$ä4��#W?	;H��T$&Yi�_`���'<k/ŗo
"�_0�x��@��<`Y�e/�7G�B��;�/�̷#F���j.Y2h�������6�W͏���ql�k�3�"ޚ��*�)n=�hf�����mI�}ڷ�I ��~���t��������O���������b>N6�֮Yhz�9��vY��9�"�6���7S�'���b�K��C��Ta��魍��=�q����J��h��A�?�5��X�z�,�BH/�^�qD���q�c������C�^�U��Wm���|]�4PGl �hF8����n耒}�i�Lo���G�=4�6ؘ��I��lnT��oG�d��4�oE|LA��Ӵ���.�i��2��(M���ֺGQ4��Ҡ(�eyRo~5a�?˿���0^��\n�+HJwW��_R�Z9`"2ob/���$y
9,�,2~��OnO�m�X��PY����7��Xg�RR7-�n5|���-��_hp�"Y.������L��IQ	()�?s$
M+iL.�_]@���Z�֬Q��u�>%.��4-]���&:(��T�6��T��xY='�S���OP���{�7�ǥ��vV����j8���97t/�hyς*��8��5�m�h�����E4��d���c��h�ѹV|*����G
�w!�$�͗�Õ�{���YX�Vp��&�
�pe-�PDs0p������O6cIp D�R.�(dN��i� ����J�����*S�����!-��䬸1�x�f$��@�mP�<j����%`%(e3}so���������d��<^[�S�N�q�(�:�`N�E�� /�T���/Q#�Fd��G��vա�_K!��T}i�bџ���������ة�y'�
�~r����d5�%��e��F|z^&u����Y����@�ި������YKk�i�6?͙q�x�]�/^S�`��0[
L�/�����* SS�¡�����%^՛6�\F����͗�1�CÂ�(ɦ������%���O�\0�v�A�R�����ӿtc�S1U��P�o���&�r��(PF��*>i�շ��!ۘO���+
�9��ח����
:$�mM�̡���_&��-$`R�f��k]7j_�\�5Ñ1�g������R��[	�gۥ�q	V��ϡYq�!H�9؟P%��2y�Y���~ȺY��OW�vX�xBG��|-T�tY�;���G�l�q��O$�թ��l���Ӝ�l��C{���'�ԢeK�9���f�
x��OAa��Ѝ���)�/X ���4�?H�eJ�r��������� b�#�9��A�[mW>w+1E��u��;��g^�
�q�\��{9����������|���M�' ƛ̈́�u��񞰣Q�^Y���c�b)�Dě�p��E�9ju�GsE�=�B�S~��Wى\�l������m�Հ�HG�In��,!k�f�b�#�v�cӒ}�� m��ju {Vw]z�/qu�NN��&����ZE��O�?���� v��-�k�mC|Y����[�G儙�e
m�f�+��� ��X�N�$������I^A�ӊ76JJX���'�������~�`��G|+�DC�8n��8����Ֆܦ�,N��秒��M�Mw�(�������=�3��-��g{���{��ʞ��bhʤFj�y����r4��obAhf���/��ux]��(�����<Js�]}�2�WQ2r���`#�a�HK���-�^�Z\dpԽS��k�?1�
2ϫ���lu���a���v	6#�C�{���3w֚�Tª�}�j��4�.E5�u��y^� ~FjlĎh�L��n�ΞI" ��,�^�ǥ�]n��d-6�F�~�$����xX�=�^e�dI![4k�3�&(#���πIv�8�Q��:�)->��T�-�Z�h�d{ZFq��T�M����J���je--"��Kk�OB%l����u�N��`�s�$��YKy���Jz��j�R�S�WU���TQ�)��9�S�ߊ��H�3�����f�P��IS~����"	��h��@�o�|�u�_کljj�h)`=�Y�w�}���^��|
 	�^�|G�ȍ}�݌��m�z��]>�D$�����\�СN�ͪ����'_�q�?y�vE䓁DV�6���K��vYHk�ݗl�"'��+	���hgE<%H�F��p�a��}/���ɷY��7��-���������V�����e�����w�{����������M/��?z���j�{;���¯K���&ce����[����s���)�+T��G5�� ռ/<�8���u�T�a�U���g��5=�zWQ��s��Z�9�XH���΃�z�\	�=�\q#��it�^��=a�H��_H�j�1���n�s��(�2��O���B��i3���iT$n��G��л�hʟ8Dl�l�sq/���.���t�U!}ι/.�M�|���2��L�R1���6$b]��vN��Aǅ��S|�4�� ���
�� �=���H���v���[���b̕���1����~^Q���N> p��F6!�x���җ�:�L�r��ԟGȽ�ԩ�R3�� �`��8 �0�nz��;��6@�Z)��NR�m;QNf��~,�ޖ��ھ�dY_x��B���sDD=��W�5�t��D`�u=��I���;_�E	�,���ܚHk�8���ӗ�/�4Z�ih���齌'G�.��PH-.���M~���]hl*z�_s�]kR����O�ݞ�>�L�#�I�k&�-+#b
�}�����Cٔp�5eZ?k����5�׆{��[C{���i-�ʶ���as׷���V����kYJBε(��g�J�DFPo  G/=<jꙋ[��=a�.!���H���;E+��=�WKL��٣����Bo���Vu"��nq)�4t,)L�#Q]W(��ks�8��Ӹ���z���i�2��&�4 �e�E"@�ϝ^T��y�#7���D�<;���ˮ�Q�`;���K�`3l�^��<��̉Y^�s�w���A��k��%_�=�a +��o��%<��Wh/���LE�����
>�o�xE{4�t'h��1/��Z����R!���LY�
<��_4&����2{O�y���x���+��Wl���G[�d����kA����$�]UX�+�%���^��H&��D_��E�Ć9��2�E��qHcu�]��xT�"hY�i���s�ՀvL�It����f`jʟ�r��5|�uN.[�����.!0���Gy�ܡ+вE���A�����;,�!�^�7e�b
yI0em�]5����qU���E/��Iy�R�t|�{̣A��pW8Q~tt� 3�{+!�T�0Ǚ-ݯ	W^�G���<�0\A1_���/��1��})��eNqFb��9���jo��
���p���#:oKO-}���>��76�-8G��͹� ������w�$�
by��L�]݆��g<M����A��o�4E�)S�q�&2bx9	�y����w���0&0�3`X�r�u���H�V L������U�֔�9��)$�6��qSKKIL ¯���C�ʵꯛ������� �@^Ycy^��9��F���Nq}@�_�ܹ,�	ڽ�x�����K}�r��;���qdFF�Ѽ�����( �*�aYZ�$�|�G���%��j����#��'�(�<�O������yq���N*�%hմ�[`�n�番���|�y����G��¡�ЕX�omr��������OH�=WH��v�d������aA��aQ<l�Op�N^zn����n<1����2�?.���|�!�C��N�gi.�m�XF2O�
���+��Z�xA/H��s��҇������v��Q�^��=�5���r�g;c�*���o�	���X����~+���P���C0�-x�@"�籶�͟WD�	^hu0�^w�kV�M*!0c@k� Z���������S�(�q9>�UͿg�Q��O�M��(��cm���.�wy������F5?��`���|�f� �,<�� 6՚:�=�'�2hn��'B��[9�$tRy�NW!��t���8�:�|B����` �^,Qߐ�;����ѣ�F����3��]��ʡ��C��D��c䈙�[�톿u��xA�#ALK�;��Ñu:�à\�Q�N�����j��U�P�g��a��;crON�d��K,+^�,���p�b����.n�z
f��I��E�y����a�U;8!�N�H�o9�����X��ёF�w1��Å^c�Pe�Cg��G���R�^�����n`�L{��!3Z��P����K��lT?HU��^Z-�Z�E(���wg�Y��@Ҝf+�����A���0OBQ�
`RI��2G�����n<��R��G[Ӵ��6��>�c���
3���R)�%�
��C��J݇�R�3����'o\S����0�-?:fw{�q�ס6s�ς[A�,~�K�����NN�!鎓7�L=p�4�"Z�j�A&�˟A�/���fW1�4�v�O��]�d�<���ݧ���xm:���9��^o~�X����*l����,K��v�z�`4������H�j_��`��\����#���m��Z����r����@�,[�PD�S������G�O�/�.+�䀤{��@�j�^�iW�N��n�MY�UN�Eƣ��'����|�m;9�A�c���q��d�ۆ������^mx�V���4b��'��O/��O<�������x��<�n>�]t�L���<�Z��G��-��j���S��_m�x����W�^��E�t<�'���ł4Bz�z�-Ɗ���~Pы��}�P�!1sO��-h����վ�WA����wz�xk9ˋ5����-��
��=���2#�r:�H� ��C�SȎΘ]w��c�$�T�����-����2b�#�O�_I�d�Ҡ,�O0Ζ��;/סLb�ō~���~Do7��x�R�ٸ4	�ͩ�0	И�!k/xD�Rb{��Ίm 3U�E>۶H5�Gm~����9@i��G���� u�͋�� �����侂
�_ BA��ohƜ��.�9P�v���B���a!���h��E4-w<	6�����F�V/�r:�?{x�Z>�a�t4��Bs�c�%e�*ww}����y�*>�C���YsJ��?�\9�5��"���ʺ���姀�]���7T��w���?�s��`2���U���V7Hhf��<�VΘ�:�����!�n:��^��n�Np��9c.���Ϸ1 �2�X0�7�7�Ь�XJ�}�Q�Y5�χ��[�T�jܥ����U����_�ks��k�?C��pDGWF�5�T�*���[�!eF�0T��{����� L�����ހHDkd��u�s���s�o�PbQ%C�2�}��O�����/��,.XHc�+��������_�p�z����70rR>�W��I��p��p�/�C�3ه�)2Qv�f~�9�ɭ��#���83�2�
��3~��D/N�*s��e
�����a�/h��@T���mg���wڄ%X߹������(@��L��`�5B�z�%	���KG�E�|�$q[F,vZFCdF&H����l߅ �;7=�l�\/T ��PЎQ	�{m��@JV�w��"G�p�ۮ��]Z��j|�W��ъ'��m (��]�G;H��2����D$hj�>����Eܗ=����+�/L<f�ct��T�D�GlW�ѕA����ס���Ն��!��E�&_lKF�u|G��8j�|˖X�Zt��&yGE�Q�G���yB�n���l�@�nބ��O�[v�hP+�E��)�I�D���a�g譂G�=S�xE�}�&�H3��J%�O��*���]��\k�Y�o��6np&͟@�\?*L�&�)8���E�RG����a�2X�>/(��2:�	)��|G>o3;	z���8�KlvF?�A�T�k���/���jI܏�]���x��p�׼Z3����U��<�M|#�~�mV�.��	{`�쮊�iӇh!K9�����y�X���%�Ϛ��+�1g�5!%2�,S��s�Kd�_c_��>OHK�:6����`v����|�h�F�e}�����}�횙88�"q����zw���Gd����g��	!�p�"��w��"��@k�(��p�m�=::�=j�'"�^�M<M��\\�����&i�"v�K�̌g�`x6��l���*+2+ƾ�͘ʵ����l���^W[݈/#+z^��dN*�/�1.�M����?(����l��DD�i9��I��j~r��.D���!n�#�N>�����P�o�nTC�n��1�k���WPU�OI�z��x�F����U/�c��/��	<ÍT��ւN`��{���2�=_�������^���<(G缈s\.wN�zw����L/5�i��5:����V/dΙ(�ƈXo?�1q�o�=;�����6��=���j��������r[',���-�c��'w��9��_05
m4�'�D�է��6��6v�U:�!���K��Пջ
*[��q,�3��0��*D�q~����V�QU`� ��\z5sD�0i���t�ș��������M��uj<d�Z�d���]rL>>�:j���0��(V�/,��ܥJ�yc#BM*�MA�#'��+�;0�6���[��l$`u1Jdz��2���d'��T����3��~�3�9Ӻ�޲M{��;y������:�C��%����6y0US�H}P��9S����m�����������L��c�贛���n�r��~�j���u7d_(�Τuq8R�c�[J7�#����+0���S�K�ĒtG��@7��K;k��Θ�Kjxc2�sQ�^=^3��q �4���e�-�>����/{�<��H��<�؊��q<Czg�H��9�2?��m�E#�R)�V=qN����T�4#���|�m�M���2�׳f��u�Xr�ַ�F��Q�Ƥٺ%�?^N���[�鄓�^��"�w��^���{R��P�mi?b���"f��+W,TR�M�-Iyko��#8�q�ܓ�{X,�g2�cE�O��ԥ�����hl�,$���*8l�[����~�B+��h�����ᖖh�#�Ass��Åjd9Z���\�VyTN����Ok$�ǎ�?��hd@��6�c%��%�K��cKS4g��M���_��x�AM�������y%%U
o��~yw����'בy���p�jF�����-b����毗=1��%ԟ��4�k����sJg�X��i������ͷ��@\���e�����Eh{(��/�X�9%�#a�a��i5Aɗ{.�M[���U����4���gB�O>[	�t���\�
�4��r ԑb}ހd��o�2����g�Ś�u1��ؗ��$B̜WI��.��
�u�2�<��E�tw�������XonX���Pe��a?vB��k��2����\��ꡃѪ]���<-�6]�8e߿�-ʺ	6&N�[��q
ۃS�b 鋅~K��bޢ�=�> �ݵ�Z���~JD�KjjAG��{��6�|�d�i�*p{���g��
h�E�_�a頬�/�2�(vl��������߾��X�:�W�r���ү�^k)���H(��bu��k��5je�Z�\e�zsX�,e�O�nѣz�}dݼ����4�1|��t�ǩ��~B�&u|���/��_��J��,��~W�6�՘�M	*TP�W��Hw~��%T�FDw�#gt�� =F�כ*�>��2�l�_o�F� ���~��ʏX���w�I�����SA�
���u\�����}��hB���˶�sh/�	������kF,CpT���9���xB��� e��X-��r3�go*z�nN�Kq�)�ѧ�}� �?Oܳ�Nu�`d����u��J?��!�eaz=VnPQ0(������i7?@�!���%noJ�܌��e�yk(:��`\���9�d���r��-�����i�.eޘ���	THS��qx�kX�����2�im$�LƦLý!��ݙ
hm4�G�r�X�>��TJ�k�.�l^���D������Q�2W����nN1�wj��ё�]�>2-^1|�l��W���$Z��6RP�8戮��Y�
��2���Zǉ_�I��8�b�s�|�yj�~.�	<wH�SڱϞxd_�9we�A�9@�9�$찑�ʤ ~uA�:��V�����.[��Ꞔ������Q�4u���gXt��`�uE�|�v�sy�>��l��NNaBT9훾Xf]j�h���dߛ�J�%W�LoYq�QL��6����M��V��7��O/܇�R�9�6�B��#�)`ErL~B�ґ^8rێ:�̿e�5���Gͤ��u�h�*.�6
y�V_t�P�TG��Y73w�����hM5���2|H��$�Q��W 56���t��ڀ�jȔ�,RY�J_q�����1�즿�����l�ighZ��H139�`�����ԈVQ'SYq�h��5Nn����k���e��Aj��ҳ���)�����p���[Z_��p:��Sų�a?�w�@!xѯ�~x@�xA'vw[��f}�Z�W��6�2��=��5*����TIpn/��_8I���ZI��LiPJ[y-�����x��|W��\���\�H|�KD�9��yc�+g�t�� J��Zv�V؆qW��y����-�{N��5���B����N�{Y����a��>��=�����l�^�R�� WS�����Z��a'�"Y�U�����Un"G����5V(\��0*"��{h���[�^�ֳ`ꜫ��'S�/PCy)<W�9�O��
��p���!z �8<�A.�q%>�D	2U�H�{_/ �������1��uU|7�H���W������][CD��������_X�~ӽ(���VL���hڹo;��t��%bs��ْɚ/��{�8��?�y�׷��2=�`��r����, ���M�'R姹�;����O*�2�K�5�����T����bSM����o#��[5����3qɌΉ��j�-�-�9��ֹ9P�Ef�BMҧ5�����hfJ�?&�p��ï0j@_�&�=�˺z�\	�U�����i�b���)=͍��<�a����ӆ�&fyw��<�������:�j[�8��%
�W�aJi�}�]W"S�/�#I{�1�w
���H��i�#X�36(Q��5�g��;��MS��S�.��[�i��^�17>�*�W�q�pz��'���2����O�J��򴴟��9���߯��W��1Rp�_~�e��Y�/����b�/UUq�<V[r��~�J�]|�A�7�����r��s��x��w W2v�N�OZ�������"H�#c��9^����'ph{��`�u�2pk��s����v��*[L�|h����C?��S�.��
���Jf�L����L�w����1��_�\e�t���Y�XU&�pkA�O��;))8��)(i�LBg>ǟ��*v(CE�Ӈ�P%��i�F��⁁�v0Bvyy��� V(/"@���v6����q��;"3�J椗�F>,�M�SغQ�c��3�dӈ��a��9��x�}!�0�镣��C�"9%/L�n@�+�!Z�s�È�Ǿĭ4n�}R�c���Q��ĥ���ޗp�R���Αډ��J����X�P�N
��B������m��<�>��:ZZDttt2}ԟ��nz�2��Ne�|��'Wn$�%�勑%'ߋȫvg��,c�'�!�n:�,^���X����r�)�I(,q����b꩏ÞT���������[_)"�":ucߣP��E����B�دǐ�6G��ˇ��N-�l�*�I�E8;;OJ�S��8����������y�?�����)�Y02�P�]�
�����u���1B^��m��}��k�NWz.E�:j�~m��@^>+s[uS�oii���D�z��p�̈V��r��VY������w6��i-:F.�"���@ծ04��!�@e�W��%������*��6��M����3�?���~�z��rC�|�<zws˖.���N�]�}$���X�sCt@�n�@�y��� �����ku���_��]q@�E����!Q��6�k��s¤|�B�*y����~^�R�'�/OmΘK���
u��*�z�I��J��r���F#���>K�|8�b�/�����f�����C>~�dSW�8�ع���N������5�9�:j�_L�l6��RB����k,������[�x͚ۏ��`��9\'ؿ�jT@���ԴM�D�rʄ����^��mM�\�VL�w˖:�59s�'�C,���U\��7�?������ZX��\(��{b�DYT	�^�6��5�=���Xu,���%�ԉ�2)(������ɥ��*�i\4df���'��<<�(4$y,E	O��Ж�@�7A����z>���M��ү�*ӷ�aG31o��z����� �u>P�gh�0A)?�P��<:�'.���'��˻_�vf�� MG?`r�%�ٲ�ܔ�ebL���I�rJz����!�g�_$}M�s$� S�:�u>3��ψ	���<�qo���+�5m��4�{c$,��861��|���)򠸵�g���p����C���Tܾ"��1Q�J��B݋���R�+��װ��C<?�_C� 3���%���է�:�v��I��ݻ��0&���R)_����@�I~3�pN�r��2�n��Q����VR�#B,2�������WZ:M`���g�+j�NtT���p�3??����ۿ�Y�Ͳ�S������(�Rso�h�2��}��x���\��B�%���~�o8ѿ�s�F�o�o0p�8��DP�K�;'ocJ��lҶD�p#à1ݱ����s����5��\tt0a2�hȄ�8��y���eT2�,����A�P.�C8�I&J����j9:j�{�@g[8�����Wg�a��֛@-"gg��.�T��H��a��s�h����,+�,w=i��>��v����� �`�w��{aCn�|�>��!X$��j�R�^_�e~inn>�f?�0�=�Z1���$�[ɸh[6
��jP��@�����S4��):^,��5������T�[�(8f�:&�4:o��ɜ�G�������8��l���������\�j������󆝰�A�L�?U'bu�!�>��H���)-�7J^mo�S�0�n;��8����F������׏�������3���S@�����HS����b���2�r'�V���69�����ʯ����խ��4��,�lI��0�q;����e��,#��v��z�ؚ���U=���VH�1��>�JBӨ�E9"�1���O�1uj��ɛ�^��ĉn:� `v�|di���(|�������'_�o͔� �T�|e�@{�LY)oI=����B͹NN�u���ޒ�������4��w<���������������2�@�I�+!T�������C�w���=���ze�h2#�X��,�F�݅�-���Q�.��D��H�ׯ7��m���7�/��eS�L�,����]��/(��� �|�|�E���+�w�J��������v������P�<���_�]�~�/��s��5��x�7m:i�P�P��\Z~s`�#`��F�N6��c9<�nn0�%�ܑ?�{ak��Q{��_�*:�9���m�X4$e̚�H5��fHf��g�ΘŲ`�U�-�.`�!�v�ɓ�Ց=�����������޵���AB��E������������_�ޟll���)jhh,,����bL�b�X�:����8�u���@�^�e>�-sj_�g�.��cR��:���Z_?��,i|Y:{��?�������6��6~�`P�7W'j��hGZ��
�����;ao����B�_bW�����������v+���������k�p�,fo&��aї9�����%. ?����c[�-m��Fc�;��_�[މ��X;�R�����"�R�~���K���������}mov��v`s�@�J��9��oo��.����9��ʜ�>�"u�B���+�J6!u�+�w+����W�Sȷp>�<�JP��x
[��;�jK���Z���2(���}�$V��S���)��f~��^�n����ɸ���3�=��bQ�^��>�qb�� �bjF۫P D�k�6��kZ�<
ٕ.D�5cvC=�����d�/"�}Y�����[Qɔ8͆88�r�XI���U|&�2�1,�RP�����
�>��i>�#E.��؀���z�ʧM�U�~.��K;)RJ���1����b�ڏ,���qνec\�c���n���P3&�1�Ҝ���\�2�j�%pJb_�u�{M@�ʔ*�������4Y=�<�?��4���y	b��5�������H�<�p�|H�s�|��v��D�wvt��� �j�ϴ�f�� ?�_ҲI`��U,q����﬌R�UN����?�o�s�|"T�C�i�\Y�w	��V�81�n&Bٔ2��5�6��	R��9��Ÿ@����`��G��5��ŵ1`#�d��h�K{Z�fA����V�Dr`ܙ��c�T����OJc����a4�Xm�fƽ�r9��y�*>́+����g�&�g�uǳ���#+i&&YǃqcUs�@��S�\�"U�s���7���&[r�o���@� � p�2�/�ӛZ��������h��/�"��վ�M�ٍ�@�r0y|D�۽r[2Lv-rQP��#G.YQ�������ߺ� "�s���o5c6��~�"A�O��Ȧ�qQ�������tqU�_SJg���PsF]C��I>�k=�2L�D��0��K�'�b+3׃�\�nT������P��-n�7�b����E"[�(2�Rc�K/w�?K���c8L��@�����}4�8�e����3Hz}�+�֭!�� ��Ds�����©;z;��SĠ(f�`�]+WlƎ��H��G0�
T;Rm�hr� �g薉d����0����K0�蘧�$J�:�@4o�bnC��?K0U�FoV���M��@����~�9#M�?��̄Eβ����'|l��M����	w�9����{� ̰���OJN�����$1]�THg�)U
�?7�6p;W6�F����`�+b�g�r�ǭ-aeUȏ����KWg�!Xh*�fy+�&���|���{3ڹ�zΥ�*B6����4*ս���k��'����	�˅��/�BeN�fҿ�ɣ�3�4H�D�Y�| u����$M� �������wk��]����$G`g�����0�(F��Px��p���@n�>TaÖ3�P/��ɡ�d�^���6�����_ƕ�_y���G�3��� r�C��,|ϛ��w	��b8YI�Z
$"Q��'^7�X�s��Cy�	.�,��)ۭ�m�Y�$ޤ���'�(��]v��=��\��?�x�h���b�osSKwR�[z��$�������������Q]��sZ�^�E&�<��=c3E���ʟ�&��~��o+�ZZ�39�[�6r
�tDD�>���oֵvE:�y+bf5����}^}�a������/7g9�ƕA��n|O�|90����r3ʈ"��ϝ�CP�՘��q�3��w�y�F�՗�x9M?��v�6H�O��N���Z^�Ϙ0��*+%�Z�`*��K���P<�C�:�7.�;��lĤ�Y�Om��1�O���ED0�N{=�m,��u��k�7�ρ;��__���
p�#!�t�����Q#�2㖘�C��"{����_���JO�u{�9x�ɤ�a�����W ��5����Cp�Cp������ݗ���K�]���	�o7��^=��������眾�}�)���<-V���C�p�R�0��`3����g@��g�,"��/�H8�����$�J������(���He�Y�nv�"\�8e��,{e�5d{����7�I���
4�n��@�����Z���w�sҺ���_�؄���I�һa��I���5�l@:������?�6����I6�߄O�����.R���7��fbS~-�f`C���do����k%t�DR�0y�f�r���@\H}�N�KB|�rv`n3N.)��gf�q�˰S"�;��?�.Z���#��r?gB��:�.��_���w~�*!Ŗ+^r���l4B�{��0�Q�Bݞ�Ľ��m����gƯ��b��w�|̇3W�Rm�9n�lW>�F�!*�w�&~��}�ڨX����f� ���h�q��?T`�LOǇ�e<[����o7�LW.�����������nñ�*lL�Ӳ�˽��Ł�/	�p6��p`��z&�7����y��k	�E� �A�<�FƟ$�Hї ��(��+��B��B{�!�ş�33A�ӵN/���)���%Z9 � �5���iݘ����R��kU��I!��Uӳ 27-Y�����5��KO���ޚ��\�UV���׋�#�3����J<��3w��Y�+2p�#��%Pr�5�چ!��vKO|�8��֧�6l�;�ZlF�Tr���fI�	[�B&g��!^FW{��d��罐R\s@噬C��뗆Dga�:I)�,j��)	��;'������rw~��+d��g:�(�1�����7l�|?���jo����cc�ǹ/�J����r=�w5�%�N�DW�nȺ�������PY�7(7SGkʡ�l�c���K	a;�!�`S1hw��m�*c�0ºI�J:\i�u$g�x�E�Z� �r2�#^]HwUgQ|:���!e�Z�p�3��q`Rc
�3pV���)^X�рb����f��?f
z���ڎ�5��w��*����8q��u���m��Ib$�niiD; p�]՗���|t� Ff[-ߖ�lX��4����?���CY['���>:��ӵa�@Q�_.�35y���B���g�L�(log���oJ��{�w̨w�$*��ʐ�n�PW4)IV�f�V����_'w[�����m,��V�>�p�l����D���J:R���W���7�B<$v�/b;�>���~���Х}��W���o#���5j�/��N��Q�2\�`Zx�����r �'Ț��AN)4> S۰����YfYa��MRc��t�ZbTV�S�}�h}�a(�e�~ȡ���)����ř?�CU��!a�8��H�,�]��2�֨�����qa�9���K2�D�m�:�t/R3ݛe����"��:m`����
��_-�g���Y$�����Α��bv��R7;>uc��� �7@����U\k�>��ў8���Z�;ߴIh�r�%���A������-?L���;j,/,�V�E�'��ӕܨ2=~��h'+��g�Nl�?l��>�7�ܱ��W�P�DCC��;B�<��r�����4��hDJ���>1_~�5hM�]k`-H�m�΁�	��VS��cI(���	�� ��I�f��W^���)��G�_J���g�ڽy|������� t�z"I���{�����p�����I��t%D+���ҡ����O�}�7�o8���A#iK�6�C���*�\��&���吖����Ď$�����OeC�O���|au��sc�\)�a,OGL����m4_W	9�,�ޥQ����Bj�r}��e�"Q��;(��o-���|+��Z�c�����%��O��YX�Z|?97X�t�a�}�>1u���R�xk~�4�ޔ��)t`�Y}JCy���X4#�k���i��_�Y��0R��e�״�4��Z�!J$/���6�L+��n�:�o6 VB��!�(J�P�Ł��)ѿ�:��ąg�`���Q�"�0��G+Ni�h�zl�S�!�%Ov���5,��ŊC��P*��uo��]�<���!�Ǘ8�V�����6#��]]K����c ���Ku�^�'��ٙ�n������^�R�ꏇ���3�%��E�tv�B�Yr>��Q�Br��
x�`��9ܪd=��JTdHj�/��c�������v��t�P��ׁ�u�۱���!o��eN��--5��V�[zMw��QS����K�w,���I�O�IO��_�W1XN�K��t�^�U�Ώֽ���*�]������L����b#c�����v�fyb��ٟ�2�:�4���f����X�=Z�������@
�,������(#�]��c�^`�zR��`����7���QL8�U\PŷN��!n���O*��Y�>�}H��z�I*��=< �����-?k��$��x�/����]���O���s6�J���L?E���8��
���? ����wƺ�cO�5��gLNB0��,(���	�ׯJ9H'�i�w��0�#�>.�#�%Hn�n����|Oօ����#��啿�/�����~�k�X�>����z�����h�<:r5��ǩ����~�h���+N��+��ǘ�!�qcI�:܉䤏�a�4	����V�4c���C�;�G����y�!���X��y��{g��<���|k�U����A���,����ȞVD��s#��A~�,������>�j/�\��Y���2��OtG�ዧ&�>Gse�{Y�NGe?��e���@	�����Uu���i�LF��v�9.�B +sVY�lR䉅N9����h�!�G?�7H�P�=L8:Y>�^-�ZW�,v��е�8S�I����깛��[�����'Bt���Fi4��כ�U92���f���Rdu�7@!Ô\ta�?�q��G��w8��<9I8ć�ꑰ�l?:IB
�=��΂QX��0�����N)t�����j����27R�-͛0�I�c��;�M����,���s�#y#�R�.�C��&��r����&������c�?]����mѽ&twE)Z�"�(�g�9mCT4P`^��h�5�/����ZM�Z��-��E?'Ӥ�^��%��dt�M��N(�|i�q&=�i�$V�fd8����_��:]�ȉ�},!��hf0Q�	�|/��S�w�ǡ%m� �@	���qxtr�ޝs�J �+Bvu�rc�*����q��[c���6$��EMY���@0�����0����/w[j�y!j�|d�r�2∌�Ƅ��F"K�DQ��_��+S����V�pF\A`��	���D���ջI�T������<`s�ͷ3�B$��w�:*#��O[҉/>�ŪYf)`֏�j�\�T~�1QQ�G�����f��o/�W��+
�p>��[��m�<k����x�L� ���)��␠�^e��C�V�u?��\�k�D��t�pe+�\�����*y0�W�c��3�������"���i�d�R�~�������+�1!ŗ�grY�K�:�BU�Q�Ws��2��G4c�N~S�L5��[��($���+��N��Q��R���m ��x��f/s�;�O\<���h���n����#��� ?���eտ�`�JPs��ԗ�tp~X?�ܰ��,c0��K0��!�� zˀK]��+JĎW�|�b�ss�2o 2ڧ/C^�](.]��Ѭ޹ɢ��ӂW���u�0=��l[��Og��wv^�8���`�Qv�؟���\`��UCzP�Ҍ��r���r�#�k��H3���9����2E��'~k�@W%�SLS�}ZᦑV"`��6ZS�u!��ߠ��*�f=�������~'�
�A�@)�k�F�}��k�{���؋f�}�H^~v��U$�ѺN��D#[A5��5�Q3��C��q��wgt�v��o9u��>��=-E�/Hg9�u���.�bش�fE.�K�!��ŀ|8-b�7�X�9�j}�˖�������"���*�EG�؅�������2L���ˆ���߆"U?�%�����ᬥ4�Q��/��rPR�qq1-�W��I�y��TxY�p�����6⚧#���l�k?��T|�nk����P`�]D�2u{���Y8D�d+a�i&k���F3D��T��'����	��.w���FB0gJ���j�
��2��.��*E��G�\��(o4�*U�z^o�>�Q�����
����O��K��6}�ڳ��9�Dl� �2��󅩹U���0½�4�Vces�5NgY����T�Z�ttML51%\�Q�nRe�KXbᛤD��x�s��'��q7G�,���t��3�ճ� ɋ�=��PB̩Z��Ω]��=՝|��ԭ��T�������Iq���!4ԙ��2d�0c�-'H�w_�M��Kc�wsh��cZA�E3(
�J�)�0J�h}����5�`#8ӑ�M��"�^�|����t�x�ǋ}��b��Qk_?������055�}��}���=��^)��y~�1�jYQ��U�P�r{����KKu:]%>���n"S��ݤ�HN�-|����1ٟB�����ܵ	��gXHG���i�|�<4
�~��u��iA�o׿�2�#���ޞDy)��t���Y��!���62D��?l��o��)�� �Ռl�ܔ�Z9!s �qZY܉�V�|��eL�u���EIw�v���姵�m���� �F�-���X`�ky��+��]UK�_��/} ����o��/��8�gEo�'�vP8��sGt�!�?�I٭^�?>!w�co�ih\v�.������9�����$��#��f�Њ�0 ��%�1'a+�*��]��"��W
����IyM]�I	9���c^�y����EE�J���������33"������~��@R,�,�۝��`��U�jD懗�h֘��9�v(�Ҽ}#?
Ӽ��#�7Uţۥq���z1�5��ֶ|��o@�	���X�ZZF���I�Y�Ʈa3ӈ�غ��o�#� �����J���n|K�O���?m/�X�����y�|��s?�x���;�aҌ8��d�S�ݭ>��Jt���,F8%p�
��=ɟK�aխ�Z����jT��`�n��r�pn��/�κG�΋���qޅ�г���3eBV,��ֻ� ѺWɝ������0c���3�����ď3|���鯛�v�W���Ъ���GCN<X���k��{q�##�4;������}�e9@T-SGI��;��?�V�Q�|���|��og�G �Q����ew���~�=/���X�hx�o�O�lT��N��ۅB��`fј�0��Pղ�Y�=�Z����^9C��t�LߙZA+
k+Ԥ��`�yY�B��[��-.<+`��D>l�e��N�<Rl7ٴ$7�<[�"�O���t�Djc)`$/�'���4I!�%,>~]�Ce;���6�QU���(X��(7��T�\!N`�U_~Q��������3c��W9��!��6���*fI�4�7�>��n��X�����>.�:|��)��������.��W���.n�w�z�|\���`�i
�|ҫ�dA�����0t	^$���_N��l�d����@^ir<�װS�E�(��4�4��9�w����s�_��:(��b"
b6/�_uUF�^\z�珮���[���A��]b	gH�.4}po��ܪ���n�}�k��m������0�5�����s"�:=�N1�6,�Ҿ�`�v�g4�y��yl�N����_!�,�s
���3͖��S�	X�۳�����5�����ι�uo��[���ƥ�՜[�Nn2��.����EV��_��C9�Ɨ��H�D�Z�LL�'o�d��nd��O�_p�w��bS�r��}R�4�7FE�e�{��Sb��ik��6�\k�.��*oC�������
�&�g��������.���N"6�G߃��jy��qk
-��fw�?(��P�� 0(�u5�k��iw�,��D�꯰Q��5<e��I,�Y��6��<z�@�A�LUM-��j{�đņ��൘e�Q^�</��\2�a-E�a_
u�&��0�B_ߏ�@x	*���3ysSy,	#RM����/�`���BKl��+\�t��
��{1�&5[$�z��ye�l�:]���2�vp$�Q�O��0�}��'��б���6Gǽ���~���ʇ����qM�o>P��F-!p�Y�W�H��`�n��'����ΐ�1���6����A0�~�H�I!N�uҨ����
�YQ�򡘜V++���UV�k��շ
�&+����� ��$�[������&��(X���U���Eu��B�IL�O�d���j�PC\XQ�j�I9|��&�l�*L��Z���n��ZN�j������
�rՖ+iH���w�6Y�a��ly�ȹr��A�8*����]���E��h:��K�H$����u��Ch���(-�]��R������D�N:��*QN��s)Rݻ���%�l(x�ߟ)��wvB��A?c�2d�do��u�::��qs�0����Ǭ�~����&�Ƅ�3�n���[0�^�:�_�IN�X/aw���y�#���Wn����f�S.�Jެ�'5�������\f���wG�'��y��q�X��oOM���Q�����,�����N=pE�Br�~�n
]b>b8�i����s~糷G�'o��b��o���^��Ja�&Y�=�k]^̾�{�@�("'��˭z"ڭ��ߚH�Ρ��ɥ�sQV�i�����q'��}�$��[���ף���TD���c�z���}p7�Y4 {BԜ��o�v��~���g�����VJ��W%��jߠg\e�Mx��)�����"�RA��< m���@J�f�A��h ��W�ZXV��(�"|F��F��B�H�9r-AD��
꓁A� �����R�>�vb ��b�(j-=����޴���}yFp��N��d��s��M[%v�ַ72DjPbON��)k�DT����,E�H��=�8^�t���?�R��� eQ.��/�eN��N"f�����2��+���E1��#���'�H轤ω,�*uJ��Y�*b��p��vu�3���Y��Gfꉽw���n�0�[#�8'vs�����}�ý�H�` ��m
l�:�S�W�.o�	ѷg"c^��4�H�D�T�d��ѕ��$��ͷ$��H;�A��������M8�4zH�K��g�m��1 _�u�{�)y$ǜP��q(k�5����l#�V����y����H�́1����V�����@��@�|�&��m�w� �����6�;��m2[0���B�5@nln&~�Ɣt!=:�-�`M�H5��16���ףF�2����]#�hƑ�iu����588���XJ�WN�w�gνʉe{���E���@ �9
�&�\MC	����PCn��r��J�j�B��j���zL�����[�(Ur���)3Wp��R���u;>Q&c(U�(�w�.F"(�{
��.SSTt�9��������^�e��P�O��Ӹs������ޞI<��#B���QZH*�j����$�
8�,öe#L�R�9�%KKP��	|?rJ̈� '�ٮxgN~��p�]�X|O\e�ǹ�p}�j�W�}���:T�QZ�%��uQ�}�(��!-Qq{/����eMǰ&�z�-]�e������8�X�ˌ�|��`�<��(�jf���^$i��#!�����Ʀ7��^�ˮ)���e�:��bBPwwt�	��7�Qv����*0��"0n�&#(L����N1]CbL����bTV�}�f�I0�}�R�0�3܊�P~�EG%��R�:x$UT�G+��ܞ�ɪ%�l�i'X���U+�,�21�Ƒw�ߖ�T�X��L��3��%I���aq�"Վ��UR������͐>:��:�t1��~���k<l�&��.h.0h��,i~��#��N�4�Ir�ΖZy�671J��A6j����H���n�4���և��}���Yjp0t�^:�i�K��&��L㧬��i���Ox̪Rh�Q �.�.|6(> W�p��hG���=C��#����@mx�5'I��>ё���9�a����ݟz���q����Y@$��p����چԣ$5��1�z�z�}#n>��i�@UC&W�RQJ`� ��#�E8�����&!���	��������	�.Q�qr
�z�{�������L7�}�?�ǂ�@@�9X
�����s�h��JgՏV��X�����M�'�#�'�9{��ju֚C�!I,,[�{s2P������Ć�U�X�̉��+���
���Oϕ/wRP�����Q�_��*8S�BS�U��b���P86��� w���$��'Ȍ{�c7����⪨XQHu��7�o����C,������J8�ǔ��?���VG5ے����0�LM���}D�?#R[k�A�'�-ނ��E�����G��72ӥQ�̇�?���Jl
cj�i�ƨ��m=����8�q��@'�[���~v��	6��n����C��p���$�ؔ��|���ӣ�����] -��ڊĞ;ؖ��l���.�HtCҸ<R�4Wa=4@*_P��Fm�Q��v&��SK�I$�zg�P^�n"����m��r <�h�"v���/�`KwBũ�ՌTfw-��wҊ)�~�߼��W+���$�+cq��ޑ|������;~����g�{��}]3۬�#h�'��w��s{���)�����8 #�R�
�t�WW��vQ9�x�¤)`��$v�mL8�{g�$![��{� X墲)�QTS�9�~��צ�`����T�lgDϏ���AF�0��
ط���k��c6�{���`�����������/���.|9J�4�r���Fb�I�Me�%:���0����r#�])��������F�{V�����âGӭ�5�V��;hk9Y��hnۦ��E��!�g�,��>�o�2��Fʯ�G�>k�:�t��Nnմ�L�[P�]��3ɸ���a�p��߮Tօ�$�q� ճh?��+i8ڟ(����$PL��G�_{�^�i2~���(��G��Hw1��S��ف�M��6�G$T����b��#$ 0�n>�+͒Z�c�:aݺߚZ�+�{�(D�u��|U��YF$HO��TEQGR�.kE*�+n�f
ڟ�t�;]��h���,ڡG!�3�\�.����dn���;�<�֫	�:�'��}q��߼<a	�Ka AQq}5|�&ܰ)M��H��DݻS[A� �:���Y塕&�/���̀�o�������?�Z#�W�ۍ���|�����eO���?�$r�M:m���"R[;I���0Y�\�B'��$9Am"Q�m�'h",fԥLA�:��D�δ
e�/��� ٌ���.g;�T�q%W�OU'�O}�8��.�c�yn�����/�13y6B��CU�Xi5��#m ^�@� ��㶄����O(����J|�iWL�c�ۦ������������p����w��Nz���1�K�����E=��}jJ�ǳI+�f�P=F��ix{j�n��
��*��~V�KFІ���Z��뿺�c 7����^"(y�0�r}g�UGz`�����Nvu%�x.��a�����p{���6�>8:2>�~����8n԰��ķ�����g�5��! p���������v��Sk�z�/_AӦ�(znQ�� ��t,؄Mx�ݧV]��p��K����p�_��qҍUT�7��Fj��0XF7 lߓo]��r(�3Y_ޝ¹�n�l�(�o��چ��]�@�2Z���({rf`�2ع�[^|�'����O�וE�a7�c�K��k���@NzX�6Y��9_Z��!ߛ�:�ڙ��W�hy�$Í�y<�5������Q,������k�H��}I����DD��b������k�u�'_%$�S��P-!�G�] �WJ��~I�c�/���1=T�C���8�J�s�dℭԞҠ�v,W��<����Ϫ��e�����w���:��ᄢM�˗����s�rKI��C��Q����'	C�C�s[Z��AUϡp�Sx�S��Vh���!�.�:΃��:���-�8+�o����#�Je|�P���dl��ZH��m��� 3/�0�����m͏��y`�G�`�iz�!�KA����P�����<��"qC
��q�تP�6�'�8O.6+�t����]S��UI��XX�Γ�ڛLd.,'
j�j���E�R�t|���xN��kB7Fq������MQJ���dI�Cgc����~��k����o[5���AA��sZ�u��)���O�9�$J��P���A;��1��Tp��B&���0ݳݤ4��"�k��2�+(�&�2��Pc=�����A�	�wn������F�U��O���.YƳi��#�r(��/j�o/��r�6Y}6�Iμ�	�n����a�U�Sл��B��╨�&:�`�	 ��<kF�?ooo� (��d�J�<�lo`B�6���󆤽����g��"4<>ٰ���7���B�ͯ�v_�[-�F�|��u11s�Y�6N���B_�ⲇ������Kl&v��ˏO��F�/+0#����a�/��M��]�.6πgK1�`f�+������t��0f?�)��W���Ĝ��~+T���}k�ة��8�jB�`��2���9�N�Є<d��z�s��}�Q~+:u�5J�d���5�����-��r/�ۅJ1�\�[��0�*{>�_�M�������5�=|�i����~1���af�Br�(kX��̍��E��oѦO 8��Å���P�����Bm��(�������X�1�����������b�Ht��9�iE�\���:|�T6L-7R��_��^�,ry ��*��Y�����b���u�Щ4`n+���6j|�t5�ͦ>�6;���bz����������{m��Q&��H�z�7
8��bed������u��ԁ��l¥Kܥ^Tҷ�5�����(���	bB%�$�
�,j�3�z%v��Ln��:@���??�б��ڡ
�yP��)�ev{REG�T��a�]l`�`4�7�PzƋ�#��ԏ:�~h���df��w��~��S=	x��#�g�"ؘȖuH(#�c�P�q/�����@��3�	�c3� �q���gX|���%�6kZ�����Q��0������&	�����<dt�}t���y}�~ˆe�uy�Y�C�8]
�SΤ���_R���w8v�?!�(^�]Z5S�8V$�������[��q����!�@��Awjv9�(񕏦>R\r�P%��\�[8�mA��I*��У��K�A^_��+3�^����W���|쭟-��&x����z>��)�ŀ2�@���v!0 N����5�������C�[��J�Ou�:�o���H5���X8�Y2�'��]�L��~�{����j�Q�T)	�7����:�jXQe�K���YF�����m�+�kV�z~���tQ"2o��?�M5w��Z�.���~̞�{�H����ݎ^p�	�͇�>�$z߃���f�̓������<�@)s�/ vv�����B��8V]7������Vԯ<��D%�CA���%���X1�9�c(�՘����e�o��eLI�AnV �oʫ;4�G�.�?�Mn;�9�*�R��#�=何=<#�"�?>qpSȰ˫�j��(� &lr橡v#^�RW�]�����b�����Vح�Q��� 9d�A�����R���)6`m����Z��%kب��,
T	š��LT�(�KaCp�|�Ҵw�)t��;1�J:U�8�0<�S�R_��J�aD��o���q���:��U���)��#�4�Л#�E����E�x.��,%8u�S��7K��|�N�6fS��u\}�Ex��K�2h�ҳ��<܍%�=v�p���lli<W��u�p�
[h�"���+-a�;[%�������G�:�8
�~�n2R݋���T�Aq6�=���ȃ�?�I�|��믏�	�Y�:��%��!�fk����c�?�֐&�cf�-�5�-U%��1�d�iF�����fW�k��(�������\Y<���N(/g�[������'��W��; ����ּX����v��W��o%���<�yo��]g�V����R�Po��att��M;8 ��qEW��>h؆���r�����2m3w���C�zg9k�$U��.��6�R�f�`���~1c�E9ǌ��F��V��qKt�#j��iK�N&��Al�h��(��,��Bʝ'��^@��#�B�&&�o�?��W��jQ;D-]���8 ��N�iZԢ�w���Q�`�Fq�^Ծ����]<��3�S�����r
l�(����4f�i)��&+w���@��
2&5 m����)Rp�k+Lc|��(q�O���-B0�$����F��D�p��~^E	������x��|z��(�$db����r�F��AL�Zh������`E�v�`��.l�=*�ָ�ᐠcg�c�4��z�E4#/y�[��e��1�0cӲ}oH
�'g������N$a�p7Ζc.!�P0y��D:nѷ�SI�*j��-�G���n���|SbZ�iV�8a��P����9�CS��*rH]�~N'�>e��Nc���)�$� �`A��05��w��3�*+a�@�+̣e9�Tޓ����ͷ��8|Z�pc� ���6~�W�(�0����U碩Gg��[�875�G�c���d�8�d4��{�>���܀N�\z��a%dd�Z���~���U��$���M�_@�u�~9So]oS��7�xXS�9�8�+��~���&���zp�w����Q�TK�����Y"HN����jI=��0�e�$�P�5��U�⽙�d숾R3`'�.k��~ �����d�b�����隍-���)	{R1S��D�x��^�%&�vf3���QBN�mHD��f�HB�߲�f����b�~�1^ �abbG��@x��l��r8xAB'
k+�?{�jR��<4�R�]�zR�i������0r��F�r�ǡL�f2h.�c�A�e{HF���o�F�ϥ�=7�q�g`���H#X�hG~��0D0qC(�f_x���Cu�H����-��*D�w�D`�ٰ&���,$�@d)�7m�j�5�l�kE�4f?������Jx���{?��Sw�y{����G��s/:��2�FDA�
U�9O�}�ĩQed�~"60n���IB��cq�'o��i	SR�S���'C~������/��� '"��� O��}�CIP�Ƃg}������p�5�=ݝ:���ה��%$�H	H�=��>+�����鉌<�i���A'8�0xi��A*TT��H�g�gl��i٩������D����}�ȯ2�o��{A��+Z$0K��� <�N`����;�hӷ�K�i�Q%�)�X�v?�O�D����6�k�	�����#��w��js�
�����ӆ���a��;#=��8u�r�Ʀ��7���ɸ��5	�%�X)�	ײ��`Z��;q�RI@j�.Z����,�����y��t��}E�����|"�u(��39�>.�����&��0�X~�IX��:^����\E���E���_nnn�
rK��h��Y7�&�3f�c�����DLcV.��!�`�h6�>��h�4����?���\���v�����Y�.(hv��3	Y�0�)M,g��L�_�Z3��B��8��Uܷ<�3�+(�3^^��������:�}%�~#�n� �K|�a�gэ�@I:�T��vgSֳ���t�D����w=J���R�'X\1v��l����_�u�Ng��Cʮ�̏��}z��;(���o���7�vҶZ�� ��9���h�S�z���/p���	�gfʯvZ �f
��뻦&������=�ôQ�·��-킟y�	-N���'��}�1_����z�/��}�_�'�w0�Z��b86GGF������0��n�d���4�?��4k����k=�;XY���������8bm��0l":�ݭ���X�)�ל��-��22];�z7Fw3I�������PͬϨ
����B��G�Ui�ǩ��Y��	��F�%�K��0>�M�Z�`/�?ru���y�����Z�z����N?�f�.r��܅!J�-�5�{�Xx�[��,�G36"�|��	~~�/��6��_�xx?��W##��sarS�������$D�����2�-�]6k"P(#�f�m��[�����0�=0��{���$����R�t��&&�>���։�H ���bu���i{?ʫ�Ӥ����l�3:ZI9鵠;�z�C4����~���Qs��.�&���@��Q�l�H.�yHC��%��& D/���	��P�?���:9 ����\Y�+˜6}oɡ�j�hZ@5	���m����J�# �{��?��wJ��%2,��#(��"\.��?�>��!��]�Gт2�f
M4���%q�H£�1qˤv�U,�&d�oiP�B���Z�Y���㛀�� �����>���tY��Of��q���>55���b�� 0�P|Yh|>�@?��\�j#R�_�L�7k��W>�J�8޴R+�w����+�{xNi�xB�JaL/>|�Io5��H2vz)U����MO�P�/6�7?g�Z��� �p��p�j���)V!	Rd fFp��?����w�����2v9�mD��D`EgǚP�^|�`''�+�\�N�x�٤���~H��n�C�*���q|_sy����VFFO���v������ب%.�rFLө莽]P`z��+��M:�Ɋ�˱�P���٬������]m����6���YN,nU*X�x�ؽ��]+�(�C΀���/��~��̂�k�ݣ1���cvn��!�FQ�e���`P]��C����5A�䈓�OӦ��(���(֧VcJ�>�
��nm�esA�Q�͍rt�ŵ��	�{ew�ljW�s�<��E�G��O������EyF27���j�v�b����
���	�EL���z^_��0vG3�������~�)Dk�T*�i1FF|�K����`�01��3�Z-��4�$4�3��x���W,�l�� �V����a�g�'g;RhE�5V���뫒 y�&������*���J�g��W�y=*����X(��Oo��G���X{a!J�ƹ�F������-0�Pnl�]p�9G�r�qc���&Q�[�������p�/vHG��@ο:��zN;`s\�R$��`f&(������U��	G�|������A�����sk�dH�T�Yѳ��h����l�B'R��͖�im`2��`_\'��ʊ1��˭䀱�fŠY�>l�����ߔ���F�����(�˔1������S�#H��ͤ*T�Ȼ ����d�j~N�����S ZkX�!?'t� �[U14Lh�]413�������7z��B�X�;����X?7�����&��z��Bm.2�Wr�[�.ΒV���zz��>�@W*�G��w��g"6M�r�a�i� �e�����7e��L�Bn��D���ʩֱ|��P��:q%���щ�N1�T���q���E�)~9/��o5�pm�p�Ϟ@�%���"N�+��8�a_��^���~u���Ѻ�S.kE�x��経� �h��Q�[W���U��ce$���m#*}��ߗ����`�-��%�"m��[s=���!<�b�[�OY9�E�R�!� ,s��  bH܀��!2�1��g�������jx��a��5r�1D_5��S���j��ìL\\܍x���m������әx�7��>_����][54����gE�o�7I�5�ꉢ�Z� /k
�a=Ůڰ$?J�{�(]��&� Hz���t�Ő��*ä�KC?�'B�����(b�DjL��'��!"iS��Ϥ�'*��3�2��X�U�@�Pbc�%t�u�)�Kw#�`N���IM�ZX]���˫|y�8��9[Qx�Ho�<\���P�sڐ�1C���������f���Q��Kp��� =�/r�v�A��,�Sڑ�!w�������|Y3v�f[ږ
��rX�\�h-�S8ևs�rD:9 ;����([]����hl3��̡�����nM�p�x�zo�v>����j#�R�W]�)m9��Db��	�sN��蕚��Q<�0.&6�GN�Ȳ�Ϥ�����Y*�
fh��DkcK�y	GG6�]�999�2�1X����G�~��L��+��Zt�������щ ���I.GGG� �f�7bC�t���*D�xޤ��L���/*���dѴ���<=���BCa"8|�ӂJ��YHt����5��x���O�e>w����lcp����)b�Fp�DKf�~D|db�4P�쓍�?7��4A���P�B&�~�#a�^�q�,@��䢊�f8 \`nn���ڽ��@ӎ�U;Y�E��6׫�b���h��%�hj��Gg0��__�X9-�Z�����kT8=_����I<�j��n[�a�����>E����lQ2��h���lV��H�=���Ÿ�]	\F�p0���G��=\;�Tت^T Y����r���ݯ���&�1@�K�����}���#��]�6��&|3�]4��2q�l�k`�FE���s�yH�&\��,��:�hli�l���m��!�-���ڮa��-!��Hw�� ��t#���ҍ�]��i��Mw~��z��C��Pֹ��sE���5�F�33��R�^�&�!�ٜ���o]��*B����I���V�B�u)��d^A%z���f���Jk�D��ν�SY��B�Td�r k��쎑Q�bx*��2��`��Z��v��8��_��BY�Թ���Z�p�2_K�=���{����G���d�o+��\����a*HK��zg˾VYLѴ�nD��3�
���'��=9����oo�oDJ��y�ϳ��}Lҳ���s�YAMB��[W���4l��ݶ�(�0?����W��%f�W �"''��X�����`<4d�勥ا�Թ@��Wʋ�s�����	ּmq��Q���*�G���ŶE9�[�{0�V���_�E!�y�YD�R�A���*�J;��m��rm^)5���H��ތXd*���]}Z�ԑ�9�/}ߗ��a==33���p��Mt6�Xaަ��6��?3�U6� ����$�-Sհ�*��KE����'撴�#N!Kb�gL��j����M���0�đ�m�ȋ��Ig���#W�@��nP�'��A��q�ۙSd�;݀Á5y�X��R�f����~���|I����=��$C���_9qJ����hMԼ���d�Ywi���84$�x��'6��I~{��"M���)��d3RR�ْF���%�����Ȗr���@���a�g�?�LP^|�%����K2�����K*#ww���Q���xm���U��p��p$;��Sp�z?|c�K�|_�^�d}}Q�Y��F��2���nw���R�Pa���a�/�K"ڽ'�]�5[_����>���uCT%[F�F�ݿ���f���3�i�|���F�����&?ur(HduY���2-��X&���(,����'�C'���Hl���O��W��I�-���(E=<��AUm\BWxF+,5\��b�
�[��)�FL����uk�͇�����9Q�2������5�s5��5�:5&��'�ĒVlT9��l�/p6\0��ب�Ă���(j-�1�-��c`��Ы��y�V��;&O`���[Q�r6��M�NQh�������*���@]����j�)�J�J\�����fx�_-(�Ωm���:p��[��Nn֮��e�^ł��;�}E���]�ll5�pr�`Mm�Q�Ɲ4K����vO�Q��a��=����Op��}tq�\��%R�?4-�2��f�7�*�����b[!zhhG%�7\�8�62ߓ���L����q��:OA�����ֱ֮2�v��훹�P��(��r`�}	5�7���<I��BC�l���9�Ρ
�e��zS�E{H�\^K�Ͳ+٣��!3��aһ{Y �s��QQW���mK���9*֨���)Tb��0�{���!NsɆG�T�?��Y���$êx�-N�
��À�NHKcH�j+VN?R=�o���B�Z���ұ�鸿�\~6{#vP�o��4B�#~�+ڽ�/�ʔ�T�?-��*#����{��?b/����+%����Mvӌc`Sly�Dh���xr~>��p�gY4VvX�l������A����D��"�O����������s����
CKY�|":4�N)k5���aq�ט�v�0�R���i�_�p��z{(����°������T*��h�C���:�ۿ-Ҹ�9�x]�ǂ�1�,��_�w�{�:(�Jٯ���W1�TC��AE�܉��l��!VA���0��yo�����SR<k�����P}��d�o/!��u�H +=��r�5�Hݤj���V�|c�j��dD=Z��{��^�����K��G���S�~f馾,#LG��G�|CCJZ�1�"]�G����h=�W�����(����?�����Wl�����Y��q��8����%���$4u&��eml�>��^z��G��|��$W},���:}���ձ�9�zODA���>R��'��x��&�a�� y�0���-��}W�+�p��x��Y
�Yq�ڙ�	k��8�2{s�'�T�P;/�����ϖ<����7bF���5�Ι�fPU�wQ�g-��0���1$�u�gR(�-v���F���{sYD��U��6�hʓ�Uu9!��6lE�䲚 7�H�O�2�����[x�k�jDP����'f�������r�
�mw`�y5C�:�9�R��'K����L���
c=�\��R�O��n��N���^�&z�����7J�t�Г`�A�"�dq)|�o�Y�\M��Yt	XM�A����1ٜi��Q'otDvw�P��ʈ_Ζu#�y�.l�A���?t��!-�	d����"����KP*����w)�㜬��0�����``@�Z���5��_҅���S��Ư��ğ�\LX��H����+HR�b��
	�yA=V�XAH��pz���'������h���2�C �������L[���$*�Ac��B�Tє��J����ug4�l�(v}���y�D����1�T{����{�)��W+�����(����v�o�9j�ϖ;�����ch�`T\���.����Q�y��e~$'eP�Z���瞺�����w�bY�Q:S���
\�v%�T�sRW��g�^��GO�
 �3��Ⱦ�/��^��{dU4�#���g�z�ՈL|"qB[�7�^u�'17x�ј�dC�(]���c�cX���Th�R^���nF�v�rN)��6�q�����͝���Y�$|ߒ*o�`L����>���
X�~����j�5�	u��i�N���HY]p8�I9��?.��®�AA����k��H�P1��
��Ȁ���m˛����o��!�����h��)��tI�Ĳ"��E�6x����W��0�����G��EF����Ʌ�����s��%RQ�)!vW�&���:��-R��I�K*\�)��b�leM���sz�B�f(��,/�ײ� &�z���]��b����n؁/�l����մ|0��ڴϚ;�j�C��:����:���|�
#5�nh�������gZ�E��bU��$,��%�q4�+��F�/^�Ew ��|�B��4���uW��(�ę�ۧ��u���F�3dK|���oc7�/[$]�w���Fg�w!�v(D/�'�o�嵇��(۪+	[��$-CD�W��4]X>Y�h"v*♓;|uV�<�%��-�,�W�iJvv�5�)*��V��7�Q��'"� e) ӱn���tt���t(��ө� rc�Yϥ�����1�D7�ĉz k��v0�w{89�d������2����	+�$%�co��w1��WW,|=�����#�a�kL	
�Z�͉��@�._"xd{e�y��G߾)2�|��􇨼��Ak�c�gA~Hg0�nXs3?PjGBBB��%ةz������p�f�K������a������E>�z���\���Ѥ3�������G�)���3{nͥk��Hz{��TipDD���èV�o�l�x�`�&�M:�e�F6�u����)��Ed7��0����\#9E�X̔L�Gm�)Z]�N��3n=<*���m�1^|�U>�I��f�G�0��V�����~�}gTI6ߩ���}��ۚ��\61��<�=|=�H�0r�I��p5�2�6#FD�k���R�'͍ĵ��ROBBH������g��P��T��{?������%�GW��G�@�%/����8~�'�'ˣ0^��C����~����D���*��I��1q2��(ގ`�:��r���|i�LD��쫃���n͉V=GA>ը]~T�p�͖�dȸ47�E���� ��2�2�!8����!q������Kt�J�Ԁ�mKo�Y�*��|�O+E�`9W��yҊ@o����\䊍	���?2TeO�ДU��b��I�<���Qu�r�`
�]w��i�$��g���F|���ϔ��>E���WF���	��~�DQΤWXlPN�5
Y�A`�N�������Sa�� d��!��kj|�=n��ӻ1�|>l*�t;��H�9�1�pg#�4�r��'���ZHb�ecTmЭ�-�����M�,Z��ap\E���>�$K�~+Y��ѫ��'>(�񉶥�������I��r��L�.���$m��+��{��cΠ��ǝ6�J�����}��F�������v�N#�wz��/*%"���Y��1XIOOҬK�X��`�C�ݧ2�i4���:!���[n����h�	�؃ϒW�N��r�M�B�0ޣ�]%չ��p�`�|����8q<c�/[�P�_��ưP��~��7�u�A�#���q߃&ei�^�%?�@i��FN���������F8-�!uXS��<o_�#�>�]�cQ�E�r��������aHL�~���>_�
<������ W/��pԨ�h˴y� i�lon������꾫�Vv%�IҸR9i>�bF��G,�eפ����XE�S�������MJM[��6��%�����ֵ�X���>&sO���������3wJ������Z
����K����O��0�/TG��	Жؕ�R�D!�1+?M� M�QP}-�����,{���;<�f6�1�|Ԣ�2��C5���s���ۓ��÷�K�Bi�(*wͼ>2�_�����&8p�ս���ۨ��r��~�) svv�Ȫv뱔S㨫��΅6~�=l1�C��2��cͩ��`�vr����4��I[�Nx%���=@m�df�T�nhP��u�]��g�@z9ɵC�Rbe\��w�>�ٶ�?C)�m>X:H<�o�5c��ÌW�����ۂ��c�7���F����Gd	{�:� ��qy`x\�Ƈ�����yf�l��}s�x�{�lڥ}�}�}su�Q��KE��;�����+��������Du���f4�B�ѣ)��_M:ϩSK�2��F6s����p�dd۠Ў!��v���o�7~�H@��Gr�^�O/k��W�%L�~s��ߞ���WE�;��}_��ƴ �[W����+0�:K%4B�X6^�f�{�����#Ô	6nV%�W|}@�o�;Ψe��/#/�a���l�VE5����\���j�i��3OG�;���\6��S���j.2��u�_�/�����w��@�i�n�*Wc;��S�B��[E�X�����vwBlvw)��#&�Q�%��l���{��3{~��;�vE��۟УRNm��l��t���τ�~6,�~]c�{yA�5���؝�3���}3�՝���>����d��|�G�-
�! ��']sܪ�&��@!Ш*+��V�8����e��7vk�A�+$��F��&�H��<�mݠ�hE�W'��P	�n��ݻ˔�}UX�"�t����8�E�-���B5�M����O���g�@O_N�(P6��C�CyʥDX�y�^���
���v��!"u ����9��MOOM߷7�/7?P��G27f�F �p��Up@�sj��b���FB�h��.kEhܹ���dx;�t7<�4�����w6˞��Q��{.��Ĉ19����|\�:��E&��DL����>�=�S�p9�X3�+���8�1�ڍ���<ߞ�	~C��+D��֗�pz�$���x����ߎz�[��ټ�A:k�� pg{#��(o��6�E�CPUd��,�i`�u
zS*W��4v��_���˂���MT�&gf�ّ��X�9�3j�d�>�ܝ��l����%��	�Gy���x�6xG���혁O�q�u�ȫ[84�	�rrJ:q��Q��x@f��d�����	�$Wn����%ڎ)����S�^'�n��L��-+���:�)3�idE�!)˺n}Xn�4cM��4��di���)�	����.��� �-�ק��lv���^)�ڰ�_��$ �/�)]ۚ���VP ՐׅT�}���n0~ty5?�a�F�vye)��A&�o����N0Eq?�omoǡ| q�M��jXv!�fi�Aɟ��/��z7��&�~p����V5L���-�Fa}	�o���bɋ��18��S'�P�������k�׬��d`��*��I,�u$��<έ�]����e+��J���7�3k��J<��%r��X���p����$�e�⽢Z�6!ɉn9쬶��4]P�b�������7�h\V��q|��·=�D������x��y�ײ���;J@%�С�᭠�,ٸ���ڄN�c����9���țm�/��������N�i&w�i���`���gՖ�y��@��ƛ��á��?8��(�o5V�\5ҩI;%#㳇!��3���GF���}L<�a�q�G!��pE�'������,�D�%�I�z3Zw�hE���X�c#������0���l���#�D�:��BK3L|��!�DR��*|i*����71|��� i�VZ?�'S�Ղ�/V���� t��Y��E�ƚ��#���j$��$�V��2G��~�(g�����-�hU���Ig��������إ�C���_�)6G������o���+�-��p0��xYUx	�x�����XZk�U4@i�ڙvd�6z1�4Q�Y�����#ƐI�~���)9����o!ʭ���.)K�#4��%�_��
�w�H�/�P�,��@n�*���9������,�q������4\ ���S�©����k<x9+IˀґC���3jk���� ����pr�7��g��y�a���ݥ�o�g0�q Gd���u[Kl��*��8�,�q蔑�Q�T��ˍ\"��I;$�H���s���-A����@Ә�!��j�&��5`E���E�D�����_�)%ipp�F�!"0}"E|�3. �V����rp~_3p�C��TE%26e;[��7K����y�ڛw7IocW������C ��~v��J#V���_�W������YBV6~r�k������+����(�&K$#��-R��jNY[�pb)�r(� *�e���C^�zݲB��.�O��-T�::$ ��:������>�3�eYx�6xW��eV�������^�M:��MD��1Mp��e�7�;o/�@S�na74v%D��9����D��x*�P�L�S���l���S�~u3^M�1��Q���Կ)Q���v������sO��-��w��
�t�U[}�5�������:�kX�z#���s�{�&yj$����4b��b��ܴz�%��4�K�B�@�-Eķ���Zr�@KQ���҆��RD����N� U�y�e����z��]������}q�K=�DZ.?/9�VV�z��X&�~9�vۋ����@���0����-��^ �D��P������ɷ@O::Y��~b� �Έ<���oH�\M��HYk�� E�>w�z�"w�·k���LG.�LDL�Z>飦Me����,��|�~�!�5�a��2�- ^�o�ݿ)������������L�t�p-]�m�v��!�Bs*~x���O�PQl��CG�J(Mm�&�\��\�[���`}īt{C��	�;&�0R|�bWO����c0�htwk�PZ�T�\��P�P4��L���ח{q��'��z�њD�{��9hEXI���d��a�ex;��WM�5�`�̖�6�t�_so�j�[����H`T����ͺX�F����k)w�e>����tpѤ΄�(O�����+��]��ȴS�s$v��{�^�q+��uw�x�F�M:2R�"���S���k9x���Ǡ�z�c���%���5E�s�M����}D�n34������`$^U�4��1�(�P_��k�M/��b���!-���w'Xˢ���1�3Y�aĨf�<�p�d���c2Ǝ���"�e�`F�eI�i;��~��h7s$~��ar����e	2��I �55��v�^ <:5�:K�갔-��'AC��--r��D���
 51$� � �{�F˝��ů���s�z���t)Vn]\�����}fk��o��/pm3��VV�i܊��t;3\r��JP�W��u�dϧ���@C�԰�5r9�QNi��Z}r�k�r2��9����[���i�ZH���Ϻ�9~�n�c���c3	azϓ��B�-3og�������+�j�����>�}��g3�(�n�KoC=���ݴ�kn�a�z���V��%�w���5��|;�&����僋�$c��z�!��e�TOc�����7���G.�_Omu~���mm���B����"\�����T����-�WF`5ޤ��Q�=.���D2�~C{c�.�;���:��b�PJ�iE�g�C.�.��;�J�K<�|A��Sf|�To ��!9
r���S�A/��tI<&s�V���&���ӱ��B6]���="�g�J��<�@�iL6�iy`��M��
~m�"<,�V��f��Ygm ������M�����z`&g:
��$�����?�C����rc��ܓl���y��y�V�4�C��x^��m�|��h��1�sR���*!Uo��I5�kj" ����W_zy�	�
���v7�b�>�=�/�Du���+����T���ۿ���Ҭ��)���]����,���i�[)�_dQ�+� Z�T��ifό���ܖ�XE�����T��k,�c�ǿ�������?,k���F��C��_�5 K*���4�ˌ�RG�3.b�H2�S& X������o��
G���`a�*����0@��x˿���!�����������-�2���?�M�7S,Ny���#��춏�R��r<O���ߕ䬚���p���n�g�PR�j?"�d��v�z����HcŽ�QAR�[<�}x[�|��: Q��ܻ��x[9�Y
p%e��(�%�l�8.�G�9�0b���MQ�N�r�o�>{��D�JmLczY1��'�> ��+�7:�>��4�v˰�B���x��N7X:�I(�q���`�K�\0֏�I'�绺bخ�#���?���%n+vǏ4a�.��fS��U���?�mT�iE�$a�8�47�������N����F��;����ᴯL����Y2���߸#`��
�w_p�>>�?+���x1!��������u�l�n�3!�"46#�x*jWFW�~����X�Ku��k�1��qͿ�k��LhQ��nN6ޡ����z����a��k����P�Yo�$�I�ysZ8>8	;��o���e�ܤ�ږs�)�s�W)M�`3n��^!��	�Zi��sc���3�av}�r�k*��+H�wk[,�b[?x�6��p6�*��
E/4�����:D#�A�K������q��[-��P�n�����"P��G�����,��(Dͫ��Ȟ�i_��R�W�i֦�2���E�XD}Ʋ~��D�F6�\h���2�n<f�ޞ�9MSɪ[idj�yE�+1�N����!I��>�x��G�e��*�;���k����gQii�(�j4~�|��Ag_Q�?[.fs���a��ĳ&28�U�f�ኛOK�5?��Io�vv��R�E��o^�h)��/��d�{�k冚>�U�����63@#�1�}>J�4�/?�WS���ͮ]+�/��\���x{t�S�s�$�yB��s��"ݯau�s@��l�W6NN��n��m�⾛_�«r1H*QLp0��ba��;�z�?-�o���ƯO�f���-���?���ډ�5�hoy�9%����V{w�#"O۫�q��A*2($�c�1I�rWv�w�x�������{3V$��k�H_���_�T��?z��=ݘ�I�@2
��;�����>���&�LSSfo��i���Jo1j�#����P��S�Y�w*�����|x�'�h�+�/�+�R��~�[f_�;-��-Ҏ���������ƕ2I]��~~#m�i��v�nk%�د�m�����e����g ���fY��d�Ļپ>2����r��5K�����[.������~�%	#
)zZ�fZ{5�b�T^��V֖b��pH ���oȼ��D�X�oF�T��jxЉ!p2�^��k9ra3E���^�4Y�~2��`��{p���إ%mm�e���?��	�f������#h��f��g�~d5�Ȗ�LϏ�r՗L�����)2�N�)��񜭞�E`aD����m~�c�;�z�?�v��jf�ǝԩP�G��cW}��JƬs���dt��7*�7��`���w�J\���x�)���~N��ӓ�����M箉������˩E���GZ�>FFT �6Z�ݮ��_y�GGz�2I��f���!��� %w�b�Q�P��7pU����d��&Q�&n���`2��O@f��p�e����DC��D�5���OD�g�1�����+��SV�GG��.����8�A,��	�ۋ��[��zӫ#�:NF�RQGGGe8����:n������}�ߜ��?����e�����H���mhÜ@�[�N�_�n%�ޝ?X��NtS��D*�ȸ��o T\����� �o�Ji;�R'VUS3u��l��Wb?
b�OJ3��&~���z�L%���/f'-�0�_F��!_^7n��!�t����R.?�/�$y�fȹ=�~]�.M��U�G�SD!�أ��M;v%?��*��J �Q�QS� ��5\d��H$��]�}�:�%�?�y��-�<@x��s���c�؁��B��3j͏m���\���Z	ږʟ���l⵬k��H|�L�%�c��x�5A��}h�������ʉ:]�J��s
z�p�D~<ͺ��e��M[��:��BEaC_��Q@���P)�&���w��y���%��1��DKS��,E(��h�&���_X�{:�-y�!A����tkcD��b*��"plL~��c��Z�7�.+0���.���Bb<�Wyu��7�A�qAI?���_?���|�c$H�h�x�]��~���l�xX�Q�����B��~��Y�,� V��6�#͏^Sc��%���/�ZC���J˅��j���=��TE�(ޑ"-��z*H��,b�����y���Mz�����e�b6.H�ңdcL�^HKj²F�L�5��ƃ�]/��[M���o�O⪿7�K��9���f�X|������t)Ywi�^"}S��,��"d�uq���t��a!�Ґ�b�\i��&�M�?i��B�ܼ�m	z�Y��ۼe����!�:4�ϴ���^�d+wji�Hf����.���x:�.�tE|���-9����l^������{�v����� �����?5H~~z�^�+���?��k/��`��y��vC<�s������C�6KWVQi�1������G���J�&��h�L:ބK����-�-��I�zL�w2=��D7�/��� mtnW3��P�P3�	���7hhhvw����:ff� Uv�LP��"�25bb�q*jQˀ��V�jОF�k=���4w��~a�~���;$��+�W�aN�\�)��Ĝ|~�&�m��7Vz=���I���K;v�W�o��
7qi��Ŀ�{�͙qE��>/D���af�j�l��Z.��_����T^Pm��37`�P{C��}�������FI%T�L�m�����l�䵶v���Ա��Bc�hĎ�~`����*��@L����6�QQ��!��3H��\���5��S�P�԰l�spx��v�� ��Ll�X"���p�Im�&��������8e�	7t����v�ł�e�:�"��@������́� ���P�.��!�*�q�`yc/�Γߩ� z��A���K�B��t]��7/O���n��O��2�)�%uL��V���.R:���F"ΐ̿���|'KqS9C_�H��6Oϑz����C�J�㢉���:�o�[=������\N����a���n��k�%ԊB�r��ףݐ���o�f�v`]�$�u��Y��$�F���I� �#��H���XG��<�)5��y�@�v?�mҹ��D
�N����3���B�*�����dϧ�-�-�1ҧ3�z��9~VV��mQTU5.��q�R3Z�ˢ��UK�Q9qqT���Γ�y��V�>�k�-3k�[��1�;��n��f�g=/p��[�^m��TM
��,YO�����0k-�uE{�Q'+���@F1���ɬ]�'s�����Q(�F��`�^},���f,�V�Y�z���&ƳŌRm3�Ums��Q��,;�bn����m+N
X�f8O���8ӌ�ͳ�!Ɗ�/�:�W�ג�w��<��P�jߖ+\ﵟX��U�l%�J��n �������7���G�[��~T�\(�&�N>�u��\��S��^�Iq�£4�_#6Ȉk�W� �=ڌ��ǒ��ya�h��>��B9"��J�PL��<�	 ��2[o���^M���GCn�ċ_5
	�ksRg~U-K��_\�W	�dȶX $�y\�&h����N���Y ��n�v;o�%ux\[G ��I�瓤��N,Z�m�� A��|{_��jC��ZG�^T
���D��e.�`q%��
���h'Tk�_�"?�0�rդ�=Bd��9�m�1|}�'9jU*d����8@.��qW����?�B�kGN���u1���Px�?ؔ��0YI�{)koan^`���o�e�3ۡwW��-�~��߀� ��AG&����V`��I�.8If@��I��<���s(�◣��X��]��a�����7���P�w?~�XK�j��t�����Ω�n��93W��6ǾQ�.�۵W	���.��-V�K�-9�00����"��s��x�C���]2>�[��ͼ��)I����Q#��-A�^]������
��J�Y��ۼ�Y1�٠x_��X�,BrUDU���!�p���k���i%�H$,��=��,n'	1+�������PQCp��I]]���W3@� a��>���0n�D��ʉ,1���-��qCj�wu�^X��5�^����,��~C.��7��ú�o�A`9�g����1�}�F�%���ˏ�tZv{�$�TUy��g��?Е��7�	��E���gy�v��'�տ7��_q�AI�G11��>�͙c5�4�5������)�u��l,�"�D������b�{	�]v����Y�;�y&��{d����^�	��{��j6��*��.'9kxɊ��
8Zơ��h�`S{�m{�;
�E;��Xx�4�F���>G�Ӣh��{?p������n�^�G׾�W̯�/���p�ll��Y��'�:� ���gT���,��e+iW����f�w43��|b8�^'��N|��9!X(����Ծ[��Ӎ��܏T�yC��Z}�`���R�Gw��x�q&'YD*9�d�̥����opc�{�����ٝA��ʭs�.z��Y�r�<U�\�럇�xxF��g��n���k���o'�L�b���`��y�Z#�P���E;R��Z����aP�c�W�B��Ph}�m��>�ڝ{�!��Ɔ����6������	�޽�򪫕onli|w�⏫~g�1�3,�#FW�L�{r��tnuAr�lXʏ�M���u#���3F��~f����f��`���7��K���;�ߚ]���C����O+�z������� �8u�xc���Uc��R	�l���hW]���l��;��j_�I;<��a���I�`ʠ-�y����pں�%�q��ļ}��{�g�:;����9熪�Կ|1�A�&8_k�@�Bh\��P�V�:��{Mۯt2�iU��v�w���,��(��\Ri+��~v	�SG4�J��-`R��	�����]ն旝r��;Ocj�2W�ObG�z�Z�lh��.ɯ�P@2���׿学ԧ$M�����ۺ#s����C�F��I���NZ��6(h���6x���s�i]X��~�2Z�`U�+�,0y��5��m�l�|<�6���"N)U��H�?4����șc��u�������R�l���]�ź��ރ��б|���7��:vk��m��0�T�Q��y���&C���� (:���-K�j%�PW(�v���ۣ�jܝ�o�;�.�>	��L(�4z�x�[#�J&4�G�����ɜ��}���Pu���\��M�.�����e\K��
�Kxy��8�Ɉ]�!��q��RB�#��x�]�������s]A��'m@��`�� ����p���̿�ڭ}������(�(gk^PSg��7]~������5^e��h�(�.���JY�ݹY�zo��	q���y�s��-D� 2�R4�!K܄jz�|B�W����W>222vP"��r1ֽ�}u8��Y��Aj�������% 7�51���*毴�׶�U*�+�-_#B�eׯ#l4V4�4�_Q�s?ּ����j��g��s-����Y��=�p n�3� ��Y�I�Vz�%�Z�������^���|#A<ߩ)l�>�s��g)j�P�ܰ�����&��4?��?�r�/#S��>[�����
���5I�Z���t��������;�<r��w��#@yꎳ��w�I�K�}�T��k��>w�m7��'}�:� ���hXhYk1�כ-st�V�ش�K�XJ��ҭH��S�u��E�ZL-ϐ�=�5E�q�$�#��Kc�["|�Y�p��F+u���)���)�q]��w�x�̧J,��,>s[q�*�z�m����yI�j���r���s4詄��p�� 6*iߋ��V\R.�����0aj�	䥠�#S�Ma�(Ĥ�'���0u�h�i�i����u`1�5�ԍ9�s�.���v�C�t��v���g��t}Dd]?�T�w��]��{��@u����ZJ��}ȶ�<�Y/S��0���@[�!2�˧�7�<=��"���1�P,�%f�rHL�.���'囗�>���q��u�O$RPV��c�T����t/eQ��"�Ъ�Ҕ��ɂ�_	ǩz��1+w��,(R��L�G��,�Q��7�2���)�Mv��� ��!�'����w��O�Џ#�b�(t�r_<~��s���3Z�j���z�M�8�ֲ����.?
>�nSԫ�ok�ds	I�{���s�8���WM}���q�L�r��*�G�ƀ�"N�w����WN�M�F�JP5V��V�̃s�v�^^$�aʒ�˓�p��@�0�QL/�,�������ː�h"�[Zm��hN�ۭ7
w�{���i���թ��	�O�!�_2Վ�y����B^Z����[LٯI���W�(�]?J�ɕ�^g�v�EG�v��i>sC��[�R�Wr0Vs�ʞQD�*a�0�ı.f�a�UB����\�A(B�m�вݠ��b��|h��q��s	]QJ��HΩ�e�t���t!<�����f���`CO!��,9���oH��>�-;�[��
�eEٚ��3��5�ب��Tux��k����?`"�ݨe�.����Mb1�L#j"B��7�+?�����q2���My�w� 0����/<�4;u��>;�d�a߬x���Q>���걞fY���������J�)#ݣ�A�x�'��0�a�t�V���G����'n�����w�x�q
�ە��d#O������ߝ�m��<�"�8/�_�@��u�x��],D�����coF�=�����Le�"+^�?oD���m}C�z�W�1�K���!�@Ϻ+6l+����P(���I`?���K�ͬ��u���,q����1o��]��' ����@��3��%�U~!��B����\{`0
BW8��[o8���QmQww����a|�;PfZ�W��8�@A1������h $<���DC��<+2}���kh�N�<5����4
��d�P���H�T�]�Zq����C k�J�� ����f9��z���w�JU�t��-�~ �ӕ		�z�5(&�K�[����BP޴C�#9�L2�z�xx��BQ�{�Hg�X��� ޢ��8O��7V�d/����:���Q`g�`^�����=��A#�T��0���mՃ�!]�'b'}���U]�fީIO�s���Q�KRc����s2�U�Aʯ��}�'"��<���"#���z_o��WEb��C3�pť��M���J,)��P��XK;��Sl3f�6�J�PH+p�<�cp����{�Y�7$�u4@=ojյ��h�҂�N9!�k����ݡqzӕ�T�]�-��3��튲�T�3-j�����a�,�K�������t������KG6���X�� k���p�b6ƀ�sR�ˬ���z�V]��K��6#��ф���x�M�Y�����
�3m������Y��=�TH]���y�څ�d�2=�4�ғ��6�fD�~hWⓉ+�%�(k'�4^m�%M��D6�\a���0��	d�N�J��k͑$g�X5
�ݞ=���-�T>t��ǩ�����4��_-@�ɇ��
�Ƌ<��6� �n����G��G�B�PP���W�ܞw[�S<����q<+<5FX�H�����E|w���9��ef��!>������-Zޗǋ��n���GZ�5_�� �Ʀy��:�!�����C>�X^	�;Zx�%u	pB@��D�yi6�X.ő� 1�s�Pr~������0�?�v��-�p�c?��=����^4"#�`�0�<ã+�:����k��_���])�qb�5�O�䕆��0����hj�{iT
�{�n�1�o�;��G~�`���C���p�~����P-v|��jQ�҃�DM���@�=�1F�~�q����fw�Zw�i�[z��5)]�7��y��3N��)��E���#ꭣ����q@:�� "�ҍ�tJ��tץ�A�����N�KHww�����~�\ֺ뜽��<�̳g>��!zz8.RZFw
ؚ���=l�S�=~�ؤ���ViU�o�(��[����Z�g���65���ھ�?c����֨i�$;���K�����WDxڷ�]`�<W!i��[��o�o��9S�q;�P�0)�Wz�#��j�#���YA��$a��0b���M�{E"6���&K��Y��t/��1W�tɗ�FbU%�����)�C�,u`���
=>������o�)F��cKz�ڰ�ȶ��d�	�g \��� _�]�n��X:��J�����_�)+tc����S�ɪ����Ah�x���dg���]`��R�1�� �B�G�F�������T��0�w/U��g�|p���,
��b������`� 益��\��7S5TK��QȂ$�>����D�Z�ϻ�Q�a	>�ɳ���E�i�}��'����%fWa��,{����`w�(kDv���	�K7�Ph���޽���A�^�%��,3���6UA��Q����^p��ڞ����L�iJ�j���Ep�@~�A�%q�~�Ulls�7��u��t�T�(^���@x�Ӏ�3�:�nz��`�o�@���٩�����P�(�NM��3�\���L UpvfE�A�i�5����sVK�@��e����0��;�I���g���=We9�U ���8S�Y	��X�/5�'�V_q�p�v�L�|Z5:��s�¾;0��8x��~K�����y���Y�����]���V������?u�\����@���������6Q��w>R��\�x��\O��J�iڻz��k[���0����E��?E����W7�T�2K�F��cN"Y�C�%�\2�Y/�^����Q��UH��1s��i�?�~-z��E�{���w��*`�l�W�_����.7Kl��B��J=Ijj����|���Ǝ�ǖ�������ɘJ��@�U���N�p���d�ˉu
z-F)d�v�{��c���F?U"5�c�wZ��1~^nL��#B����(�V�T��:bOp�fdg�-�[� �0>Y��ip�l�������
���$���}P~M���*��d>��C� ��K9Vi$��\kS��6c��q�A{���&��ǜ��<�e6�މ�ы.�ĥwgV�t銲��GaFҭ��=$�i-	�+�+1��p��R�>ެ�oɟ:�8מ���F����l~t��?�}7I�����kv��p����x�4��a�|�c���{FOI��h�����%,��S�gKGr|�x�m�me���W����h��?=+��j�t�&�{f�}��B���0Qz���'*�EuI8i�f
C����0���%���j���L�>lĈ+��@�xS�'�
&|;���5Cy�9�+:>.�2z���w�=Na	�K��;PDv�9��_�E��z'������E�O!����.y)�`��B�~� R����E��ܠ���D�\�3�e��}a
l}�$��C��f �]�R����=�����ԯF0cv3R	�_&7u�]���Ven��Wp�찒�<�W��:stKR՜���C}Z��$��Wz����v?��E���_��?u�}�|9Ϛ�!��O�׶��Mnz=E�;u6���ֱ�;컨ٳB )3�S1���|�Z��ˣc8K�2i�e�k�o�&�'����ir��oS�}�lF���`�ɀ�a�2w�`�}�VR������jة�w�W�m.��a�>�o�R �;;>!�d��+Y�_$""�����F��_�P�x���P�L�-���kQQQ�k����c6²b���jf� �V�/��ퟛ}8z�j;OF��b�7�cX����������%�1���;���ВXO�A�1�mZ�������׼�1b�6�}�M�|��9��6�I��0`�>��W�BYNm�p���HE��l����i댒�Q�O��*"i�Ob��|��k�����������Pii��ь�
l��e|f��	�J�Ji
7"���|��(~(����UC����܈��������E�����e`��
��^Pцr��	�{�q| mp���m)����a>�U�t�~ӱ)�
|7VPLd���K�E�������CV�(.$w���>�U�@s��H)e���$�a*;$���N�	�%��^
�rh)Ƒ�g(�����@�����z��i?��ؘqѡ���1����֙3F_+�n�lti���]�=DCMm��I< v0}�R)�\{|���?5�4�C�qؒ.���'S<��ܘJ�N�]���cE���2F�]�s<���^W��H
FTL�\k�	���,�|��+��$� K���mi1B�ii~>�Pr�뺂�$pf��G6���A�iȬ�FJ
�T+��`�n��vzMU&")���/�\���L��#�Jd���o���<�ҷ;�!y�<D"ya�'��T�qC�&����C�bF3�����&+����S�G���~�!�/�h�H�,�$����Z��|�kz_����iX;��b��&�ƪ'E�=��x�4��eV	U.��mQ��̗�u3��K����=9m��ߔ1�Z�p
�4(��f�Y[s��`�X�h��-/\�Ea�jq�� ���4�]`�S�k�M�?f�Y#Ѵ���i<g=��%1z��|,>Vk��X�P�>�@��hAj� ���b�G�U�������ƒ�9��ׯW��.��γ�w�������Ҫ��hR���P�\BBB�����o��&&Vu����`X H���z[�]���^���}5j^��8����|��U����M�ý���8&���5�Cw�Y�8#F?7I�7.�1DXIQښn��Gy�4�]���~ge�S둌����(��"����U?��b�����9�4��&j!��nu�[V}4	�$J���_H�H́���es��8�l��<�17	TI���[[[�}PN�䢟A,�MU �K��$>��D�׳���)@��~��d��R��VY��*S��͠��2ER��Ҽ����9��\�D�u��n�̎�?A5�k+%+�/G_���K���a�/�L�c���⠳R���GU�;�ýB9I� HUW�����<'� @F�����*�������Px¥�ځ:�՗wW�<3�A'k�o3���c�̜���ol.pjFC�oC?GT�.��L��z���^�=86\�a�W�{uE&"n�X#�8��9�H߄q�5�=F��ڳ�~���]�a]�E���z����)$	��X���7P�����g6Rw(�x�\,�av���xR]�� �o��
D� ����+@�*�H�3�_��kp�˜x]�G��RӬQ��s�p�hr�{UC����AU��~��d�wKk�����m�K2��s;�o�>��|�#��6|�nUg�iv���@�'C�<���Gg���d��j�n���]M*��iϼ�apĮ��f��}�t�
Q�ZA%��b#������}��0��׹�kc��>�V]x����*�������ժ�m�ݖ^S[�K����丫� ڲ!k+8=|��*�Ę�:�9��3����H1e��$C��8�8�q��f����?��*F��پ/������ջ~��]C�����c��S}���2\Ҡ"�bSF3�5���DE���>�-��	;n4�ݭa�eV��^�n��5�V%D�9��� r�|�M��Zfw�Y�N��']�:)�+���y�Ar1���;I���E���9+ƛ��(�z�
����!a��e����n���=u���cg���jwd�ò�_�n7YЃms�{PG��G�qs��Gr�ˎW�<�ʏ�����£*�_r��Լ�ڻ���2 ��Q��Cp���!�&$H�g*���
9jW!���Լ�b��+Y�
zuU.F Lk:�<4���&����e�6��g�	�}^O�j��`*)Cc��.YQo�����2����}�OoKqh)�����۸n(�;�ջ@�~v�\gE6����Z�\��us� �����q|D[���?��Y��o��r��<ρ:��fqG����e,� �	LH�q�g��-B$����k�o�<J4:ƨ̡�nʴ5�b�!�m��ݝ,�}���e+ßBY�1�\T>)	�n�5bj�;!r�/-���t��:�^�|�����e
,g)k�{2ތ !q%�L`ECA�	y�#-�Ul��®M��̈E�V�x��
�{��u���\��jW�4ݤ4��l,>a	b�DP�j�?��v`��i�����a�^L%�;	b���Q�ӚX:��Z� �D��/�Ò�Ҷ��99��U�L���D�eK��g��܆�!��!Pk1�mX<���p7�k%jj\\0Ĳ��
�������������Y��*)Q�;�\�� ��旰�*�9�q� v}̢o��y�6l�Xv����jF������]g,��U~��V��bcq��9�iz��]�]�Tn��N�wȼ�
M�R�i�9V�s�dΦ�\/ߗ�u6��허���+��Vt� �,��%��вM�]⎻���G�[�ʹe�Iܖ`r�+�A�
?��'��[��y�<�]�B�[�ފmD�IX�-o�-����~�4���2fFO�3NOWf�5�lU/�N-*����?/�Ő��A,$H�Qp7��10���I�c�}�GQ=�Pʬ����][W�z��!��PM.������ʙXx������9ˌ���Ē�V�!妖h�nY;}��>:�â�;����d����fd���QӤgͳO��Y&GlY�-'�C��$���7�8\6�N��<WB���݀)���&&�`�l�.�D��Qf�Ƣ��OWB�d�o0*��3k�K��A:��`8Q��n��^ ǭ�� x���O%a+uZ[�*�z1.#�]{/"@�G�hĀog��n���G�OJ�������R�>F����A:_C���<o�"y��5D��5N��7M�0����c �po+��8d�����,e��X��A�yϩn�@"U��F�� ������:_���z�������<�De')����f�=�>֬�e��W�#��#i��.��Q�ߤ�Q�tϚ�l�O���T*̏L��\S�ԉ�~\�Fh;-	Iօ�c�qp��G<Ǩ����"�g��52�蝖nF��w.>�li��U�
��������9��wn�	zm\?��H������ߜ�`����O�m���|^3-��L��Fh����{��'�(6D�r��� T���s��4'��<{v��q��)�6_�e��<<_�pE�Z��7xm�z�[�m/Zq��\i�/�Z���:��ۚ���g߽�$f����F�4�1��Wթ�'��w�?��0���r�/�ǡ�b
/���ql����=�%X�ݐ����j ��|Ps�Je�#��;�Ɛ9�`2���R[�)�tm;Qo����~]�4�K�K��eA�E��F�-_���3�{ktؓ�����/W<���	g������an�De� a�n�fJ�v:����3�,�	�
��;�e�����~\p��K�a1�cyL1$& 7E��ވ��b�@/"��&Wg�D*�����t�k�}{E|]��*ŷ,r�l�\W�H��Yq��s����q#N<<<�s�~�7g[`9��tcp���B�b���氤�9ܖ/��	�TH���a+W��*��I,�a�Y���텣�KY�֣~��"���&�9��(h��#W�R�+�.��Q^c�b�H1�8��tAf2!%L���9���R���"�Y�;��+2�r�4Y<0�Wʜ�߷xP	�h����T8�����D��U���>�^��<�
>�� FTe9���*\����7	��%~���`�A��jwߨ皵gQ�tP����m��fq�,�Z��xA5X��UX���[���+�����c��>�90R�,��,�D<��u9&���ѣ!ٜ�H{Y���A�����>yzt����p��^� �c�J��� W���+�?���Y�1}���s��Ou*�����CG�y��y(\����[q����
���⦛�,��)�Ex�����I�F����x�q+Nu*L�jX	��4.��ٱ�Q��U`k_~��{��u �J�,,]��p ������ϯ|q����>�y)�k�����m�s�"ˤ}M�"�,&�;�
��,%($��y��g��,�?[NMz��3OM�8kE*�a�NI�Q'I��8�P���אE��
�&�tm��(L�
&Bg쯹�V���		6z�#��T���ޯ�")�_p����	%Ѩ��u��N�����|8��h�ݛ+��*aN�j�/wB���5Н"�r��ؤA*�O$��)�`����(` ���
*@6���}ç��y3ב�}��%is2���Y���s�����5m��9��F ���᲻�u�xj���o�EHct0���!�
�U�ڌ�
e�NL�P�r���D��=J,Q1ҳ�2P3���XA� �/�03��֗�E��!$e�9��[?w�p�0w�
 �z(Id3�� �uX_������w���3�M�nG*�d
{�Lu%ŷ�%ă�|��!��:-&�R6�/������5����LÍDF$�߬�d��k��N8���\a2��HW�m��H1��㕮_Q��j|{)��KPC�f��k6�Z'k�`�7Z�Æ-��P,�݂���#�t��$!��G˔ �_�[qo<���I�_�΀�h����;fl��Qi�&F`�PW_�ih֘�+��]����Aٽ��2ϒ#�$�F�P4�w�g\�R7�z�K[�)�8����Fv�"6Y�o&W�s-Q�l$�
��-����>o�GT��ſ���趤��L����u�N�%�S�u�~��]���N��L �V?[��:��R��s�$R����'�2�y���)�d2Э��#�'����`�N����E�*x� J����6�aར�U�s$���|8a��G
o�G3��nFS+4P�"�(Y.���Ė�C|�u��vGW*�rGS�C�ً���F�v5NY�=����t�=��
,f�R��� ���Nxv27`+�y��"��o�P�
���HǤz&�f!]'S��>ajv�$�4/��#�	,�y��[���hVP�7
>�iV�q<]�R'0e��K�$��f���w��_��FV��x��r�(Lj%����!E�/?=,�9PhY�S����;0P��������1s�=�Lv�T2�o^��h�I>p��ٲ���7��-��
Lm�h��S,�9��=��s�Iɖv�� ���jͪ��M�:s���*�B6�'y��W��o�K���p�
���$�`\i�ؗ�����A���t�>���$�v�m���������*�y?�A0��	�do	�J�>�|[���� ����}!�{���&��'�z;�$*��~֋-��hn���&��y�����>8ѻMC@� n����� ��ӁLL冞7�y���@J��3�T�ߔy��O�S��
Y���Ʈ05�J�ɀ�n�:e��qH�����:w�zp��G��w~�҄����|Gf��] {�<�U�7�45	,Fӣ��#N���2���������"g�R�ru��n��E6��m 5Q��%;h�9n,6H��fƩ�j�ۑ��v�Uճ�#�v�+�Hݓ`$�	�Ǚ7P।���vw\�Xr�-�)�=59���Ȼ9�Id�	����Z�˺�����^ as �nMIkkSrVx�x��(�y}QFo�j<ﶽA&���Ju�$S�����7����۰��A��2�/��pw_S�@=Mk^���5���2eT�}��@����:,��,�zc}��	�f�f�T/ܿ^a���r4I��|s��T��?]8~��el��S���p\hp���;�r��߰*�r6F��,e��7-�v�ڤ~�ԃ�����2�WݴZ���\_�l�/�p��-m�a��)�5�7��ؼ����F��w��j�d�U=�*��Ab���;��Z�	b�ύxÜ�~<B"�sRs_
�T�����}пhjj��3�?W^ic1��wu�^��&��S�����O���ah��ە�:��U;h�x����nFnU�e������߾�$�|��4	#���!��M.�����i���Z%�
��>O\�D޸#K�&3��t�%P���k�=M�Q�����Zѱ_܄�Bg�CC}��|��|�T ���,�F�������X��)Yn��f���`j��a���v�_غ�� lJ�� �WG_�,���� ���Y��3�TDn�t	6|ߙ�l�mْeҶ��x��G���WU/���<Q���������2@F�(��y���r�ߢ�Ҏ˳�o(4�g��!����¢%]�Ȱ�1^��1��⧟�p��)m@]�����ѵNlQ�����\=X� �8ؒ ���<R=T;��"�ˬĘHXM����5R�3��¡��@Y�i�NM޳�SZ����D��j��S��I���(��1<��C��[��v�+��"tL���
�u���F�(�m̻_z�Qc�a�^m�L.ΰԶN�~u/��,^bĂ*�4Ψ��oI�RG,�����{���Hr�dhr��u'$��p)+4�P�%��jz��9�&�S�!���XA�Ʃ��D�|��}E(#�{*e�}B�^�e)wE��ƺ9DS����)-:�/��6Q(+&��i�'"ۍ	/��
�F6
Q ̟M�a���C'T�F,�q�Igp����~�S�[��M�@x��{~�Ł�mrs��J@�g#h�CW8�O{��j��&��r��*�����ޢCó�/߀Y�{ȼd�J�qc�Oc���w�4��u*J�����n�a��!�A~�z�Qt}"Yf��;Q�PD���j��c�	��p�:z�vW��)��J�|a�=r����,���tm�E��?X�ykO��*u0ʡ�F^�<2�}bAw`�#�E�Y;5����сQ���R��g�9�}{�U4`��$��������Kv�|�:�s�$s�Χ�ۤ��Y�֣��:�ڰ+�_��gX�Q� ��T�J���I}D��᯶�9���H\�ѵƄ[�N�^+@�V3�&���ƙ���*ճܫT�f8� V�i���Ov�Z�z�t9�B�`����.LW�>'�
Ŧ|N�M��W�Ķ��>�4~ɝ�=@>��Fi'*$���c���:�w�p�%�7&j��8�(Oh���/�:18�!z�:��a<��0>�;�a�#!�WU��P�?2������r�i]���n��`��K���"������>�<5q���#x��L��f�y��A(�=���"�������P0�	��\\\�}�ƚ�p7��$�)2�r�[Ը���~a;M���B�� 9����S-��Wu�ce�s;�O��o0���kM���/l��Z��G�_Ù�K0����X̥�i��[H0��Cg�H�AN�q۷U�n\)0@ ΄�7řs��k��өw�6�9�c ���lpն�`�_�W�b�G��	��;����
�*ݑ�����Y��?'�a��Q��-��J����	?vLC+�-�_mb;a����JD|������S�a����c����ή��M{���������oiM~�H�%���"Q�Q�Y�(s��.�G�G>�)��ڶ9"�4;�>FCX�i]���2[��A�5�@�~����v�2z�2��Zc \�	+)�E�����C��of��A�b��f��)c%@��S�1+הoy̶�RrYe�������V��5����{PO&���Ʃ�E�C x�W�G-T핧��f��c�� 6z�qb��9IG��yR[�Gx&�@���<ׯ쬬�.��/)�����3�2C���������, �����	)�������\�Ww��>��Ԋ$�u��Fc���P��������u�V.�e7.��.�-����u-c�42��H��k���X�:�;� @g$R\����L�����ӭ��C����W�a��N�j^�^!Qv�V8�G���L��e�����m�x9��9��Ф�0뇆�d�P�ƈ�F��8��!V)__apѯ��)����mo�W"߸#4�(�>���]�f�����ݚZ����Y>E�
/��xӇo�� ��y���2��\�^����_�8��	���C���qK�%j�*0��P�U^f�`��n��5z��4�_}�snఞd�����乆ŢW�)�q�c���AN���33`C�X��/=.]t���.����y�����f?��LB��x�c#ݧ�z�#��������R?;�N4���Y��'��EO���%�+\wt~8���JD��~ʢRw�4F#9U��C�Vֿ=�����s����5،߆Vz0P���R1T�n1!v�6Xʈ����}فkL[�bCE �ρZ��Fvph��`����1���9(`UJ��"��W
8b�:o}���%����W6��?�H�`f�b)	&t�ϟ����P�j�&,�Y	|���+q��S*zp�kʟ��6G�Z	fA��y���+�4F	f��ψϚ+�j��|���Ls��IV,Sk��e�͎S�ڠ��s+ͣ�v��ب������Z���2�h�-- 惫dV���#�fdv�b��X��y��i�VW�J�ѯ^��c�N�p�c�2���ee4�լz(^�va�D��ED�i��Ӵt�/B�:]{V���y�eo��z8T�-�L��=G��B�@>��s3�>�љ���-�[�7�(^zv��G�x��h��,:�pg�Ý��/7�Fo�;l<�@��B��E��tw� ��Q`�7�~��l�4�4 8y:�i����2C[��V.Wٚˋǣ���o�!�� C���=6�u��#��ы������֒�)�J�]��ޘf\��"F�Q.�v�.w�2w�:�9�:[yMg5O��k�- ������L�.��B'�Ee�h �2ddc�	F�g��������z1�Ü�]��5N:����`c$��"	Wp2�k�}&�I�.&칺���6U���T�w�"�w�`y�AI:�t�[y��� H��ҽ��m�=���e�Ne�v̿����j��)�,�B6�(��&i�5���$�k̦g}�)�>�Z�%��������.��!�'�Z۹�$#?��s��do��'0p�%���;��c">EfJHs��̏�>LYJ�~�d�h�ńjIA�s���� ʬ��\�*l��3�_�K�mc�<ۤ��D��o?g�cr)m�[�!XM��\2�	d�DH�jR?'�
'i4�=`q�Ͷ�
�s�}�4��`D|��x�����}���'z�H�(���C /HĽz�q��g�¬w�~ܧh�N�k ���]��
O1�`�Ʀ����IզQ�L�c�=��X��'�{��v8�O@8��S�5�\j��Lį����!_�������'+�C[�Ow��a�'yu���Rqu���u�4D�Y� � �c
� ������1c�L��6��u���sjk	떼�K�/߃�j�Zn����|eq^�;i08bƀm��#TUT�\�����*�O�\�'I�	ͺ����c��1��r!0,���!�N���� � mD�����|�����M�g������E�������`S��v�Ě�x����E�8X�)8��łEٹU.����� c(w�RۇXYY�M�譕* �JIS����XB��k4�T'd8h��`���o~�?̸��CJ��W�_Z(E�E	���Xc���e޺yI���r�B*�?G�J���^�t�*יY�R��Z�F�V=���r�d/j-p�]��{\S���1�1�+�xNo�Mw*�"#��.H��C\\��>4T%MR��YF���R�s�Yp�:��VU�Ȓp[dVT�i�t0�56C��m�
������������y�ݻ�Vm��FmI�.ڷr~<3��d��ъ�X���B^|w/����#~��]6�U���>��qܗ��KZx2��@����c�jw���޵���{�YX̝��%b��x�i�p1?�-��^��3�Q_*��)������CJ��\.���`�w�@
������Z/�An"z���qhA�|�7Yk<�Y���q�k�|�S�ԔyUl�J��l ��M�ܲ~�ᯡ�~ĕ�����_ ��
��p @������x�Wǉ`�L ��y����(cɣ�&�+kmބݰE�8D�@ԀLƾ�o<H���pꇅ�b����$�M4����|�ڛ��3F_�I�YY�{�%�66��Η���s���opr�~�]���1�<���#�� ;"Xx������H�R�:�����F$��c�/���..z_�D���`펃(7\���VWCEL*3B88$��!~�_&� ��_�c�� ���!܄�KRYY]�g?X�����)u�p�/sZ���a�������9_E$��PL$di�K�`��é�R��U�\Cq� ���^��śƯ�5��{�F$|u�5Ҍ�NL����ӝ�:愎�%�I�DYݔ_��p�<�lŌY�������\�u;�`
ͥ��(۷��&�|�)��]f�{c9�{oBB�Z���f�:��_�٤~}�����d�F��;[a�t��
���P���r� ��	�-�9�?����=c�W:��(L͗n���մ�3�\���tG���ś`3�E,~VL �'�;gg���d<żԵv�JT4���+��u����R�>���!��#_���;;��&0���5a�����\p$���̀����<`�9�^�D��s��z�:A=��,�e�������%64�V�)S��|/�Q��x�b��`���9��5�Yi'\m�-:���U������1��］n�	l�	Zb��&�du��������dfE5��+x�Ӆ[�H�g��������(��La�u�:��=�噧����4ع�׻�����C(
6�O#Y�����bu����HD1���>=�Y���`-�������!~S����:�S�%�@��&��2E"6��Y1���5�5�ru����v$z�u7�[�rMCAa�-��2��R[Gmt튞+�z��4q��	�E$q�HM�L�O���Z���#�����T�T�~��]��;����`"x$��z��1�nُp@��ݘ��%��444���9����F��� �ɮ!����n��8���0�Uɰ�]��������h��}������U!����K6��~k�9����S�2B��e��P��£�����:U<��N������Jy�����|��-"��F*�|��"YΊ�t!���t�������*M>X�\�i�g��"�����/ɴFs����0�9��n�'+a���L	��v�t������j���񜷝���s����{6v6��oz��L0wW�^u[����S>��c��h��Y�s�����~P��Yu����9%���6�Y�l�<�g�膳.F)��i-j�Z1��eyL� ���@M*Y� �~:S丠�Q%����]
�J�R�Cӧ�0�N�l����ޡW�����E�CBB��'��g#BG�Tu_���W)��ފ���%i��
/V�^�ޅiW8οw�&'}h�"ߖ��Н�2��?n��GC�y��Jl��*�`W���v��#��ga� �C=��ټ�/H]��P����|�����^���B�W�g/�D�G}Ԩ�H^͊��L`Xg˹@��T����z)� r00��a��J|��%i�2�lx�j��E`�^{l1��}����ډ1�ܜ����YS>]�������d�z�Cp̥ d�RD;	6�a`eE��>��xF4��]=�$Ur �z���v���#��H �Y	j����^�?%��)����;����?L�K�Z�5��Ϯ��d��	����G��� i���$����WR�	:�3cp%b!}K簅��!2�g�Æ�/y�_�P��8R!?'O���F�k�����}�h�&n�������*Ҡ"���`��PJ�|y�E������ŝ="BB�'�]|%�# ���3����o���-��D�\���a��/�)�[)�كM0>hu�O_*V�ǻ�Jt�����_m!�f�Q�u���:J��NR�����\�1K��	Y���Zz�A��:��9޿`�Ͷ;� V�U5�Q�U���¤!��ώL&)�]�6��=}�X'��=m��qpWtr��4Nk=+�0�N�C+�iŬ3��AX�3��ҹ��og*DQ�h�;�=�������C C�A-�`4��*>'ܿ�p#�;�$	�M����+b��lJP#�N�������sC[�\�xv5�([K^f��%����9�Yx�F��븂_���܇Wh^T,������ld��`�3^�,%,��sٰa�����UI��pX������S���t,����H��B�H˽/���P���) ��N!���LW��0���O����i��Ɯ�>L,w�-�ʈ�p?�<EQr$nG���{ɘ�;��^mŮQ
(�X/�����+' ���M��Q�������لs�>��憎���tn��:k]�4��/���>�YEƮWI�^C�\�R��Jv$[�4�A��ݥ	�=�J��R��S���ڷ�t9$^9����c����B��G[CF3� v�T��l(.ao}4��P�G)�����J�8�u�]�����F��,�aL�<��>�{@yy-0�:%�@�P<�B������agAb�V��$*����C&�9q�YrY2W�Ϛ?^y�s����x�(@�ܑ�]���?r2��B̥3�`WOs�goD5���bs��<&�>��R�pP�2Pe�G����pG�純���.=�_kZ�^�D�@/S�Ⱦ���g�{��o��s��B���ÒBh�������֒Ȗ���@̂_:}�: -�$�A)�o�VE/E'`��Di(T��2��ϯw`KhUmm*O�������ꛜU�D�g�ӈ�t3�(<�P��r���+�D �y��b�Z �7�z2�K�+l4�@���i�+���%�+Z'��EG�f���P��o�h =��&��Y�'�ޓ��$�q��fv���2��,�	�39�ً˨�
���ٚ=�,:{a���������:�����
x9 =u�+����D�"�X"e������[ߩ���t�����n�+�p:x�wA�dy��ј��e[S�M"���8>s�Iz�&���ύq�ɳ�2�3�!�g����[+	�yN�+���xů�#�������ƻ[�(�{�^�.$��/^�_�xE��pN�f�U����+��{�z�)�M���u���S��V<�*|I
;������H���'hmO�=�r�����$�޷�ς��qO�t��J{Ӎg?x�����9����s1��0�LT}��R���~7ˍ�~��������	N��8x�2=N����<�<�p>k�)�S(-!q9#�<�׺��m�hB�c���g��*Kt�,�?��ͳ�E�Me�뤧H�M�3,�hͭ�=ؘ�,(�}�[ׄ�ܪdD���oKן��r
D��5��
5=H��Q�ӋN�[�d��N��@�����d�y�ls1v�����|��b��ڢ>�
s7�q�|�;�3Ɠ��'��i-5�$>��j����=���$t�_���l���Nͥ���b��}�1f��4/�*	��ċ��\=7_*�GXf8�bd�~9��Do����^��a�yL�����d�'�MH6�j��H;8g U&���BZ������L�O�D�zZE��{������q�G��$R�2u���Z\��Ŧ* �"!$)9ހ--8�|�z��({��b9����Ho���̍G�箳�
��)��~��fs��_[��@�t%ɷv�рQ)����	��h$WJ<+=K�C_�x�0[�j�%��<\�<�z�?�-Rͺ��]R��
�?���]��*�2�繽���m��*�)2z����+8���`=N���3�!�*�A�1l��\��8)|2ff�pвяK%u[���E�R��g���%nˡN�e6��勌��X���ݕ�8%JP�!s�|k��}���78��Y�=f�4>CI�	J��&�7э�J��P��<������4�D�Nn^5�Ҁ$�fK����"A�{�lM�/H��Ӟ�.����;;�`�*�QSX�8|��W���1�%0Yzrj�`�����"�B"�fS蟃�5�J��!r���53"}�4FV.M˅�%�`�fJ	�L1zP'�V�Sa��wVdUy.���7�0�'�Qؔo�\�bM�i'_��we���8��;two�T{�����5:�z\^=�#��=�Qs�S떔��
]#�>U~"��o��P?�]��Ib=�������m�X6���pa~�c[`#��h�&�t4_����ؐ�#)>�C/>�,r�?��/�	24Kw��� �0�d��Ƞ�
��.�&�^ҕ�PY�(�����Md�%��%y�eލ3FM#9{������ub�ux�%�!����ӹ�0��_�T������A������ظQ�Ŝfm��jv?^���f�,�^X��I,~ej��:��f]0�l�����>��-�}螝�ǒ��V�f����`e����E�Z��ʢ�k�#���b��F?q����@x��j���Wc��,]�ćüۼ�>�d���`IWt5�Ftn�y2%���[0�_�}g��h�-r��V�F�8�e){2H����*��.j�9z؂~�K�̞�����rd]�oo�"��qNξ=ݑ��I�v��~c��p���?��I)��πW��������:1�����A��5�A����������yoC��UTk�".��x�X�uf>�;#[F�k�g�v �ԕ7�?���ɰ$��t�EJ�����R�R�0B�� D	�1�Fb��ݽь�{������������u]��,r�c�-to�r`�-�+��%K��������׆nC��[ ��3JKKw�^0�e�>8	����tIC��U.iI�)0w�W�y%as����L�#O�,�,��H)6��R�sϫR*�G��;Wcuԅ��u/,�E�ȴ����Y&�;}���I��_w
w��g}u{/t�c�I�Ȁ�(���>&|`x:h�.f��Y�~w����?"l�v�qMj���.�s���R=.��p��U� �Ŝ�r*�(����;�Hoz�9�O��z_FkT�*Ro4�ғ���"�����P%��D{�l�E�A��E��" =i(o��&�ZN<`}Z���Ģ�&�����\�L遆&œ�<GE%W�e����%V�t׷o��t�/	�N�H~z�*�=�c�;��#������MлW�5{��7�����4��d�"g�O��� �3�*�t�h�+����Xzϖ����1���37�U?Z!7���.Z\H�{x�-�d����Qū��/`0���isoo�L��&��aMq�E�`uN‏����Մ��H�5ت�ŹʞF�l�h���[	�NC�(�d��P�%�~��o�$��ݽ�z���6������}��ʸ�n�\Oi�1U�5��/D���Q}X�B��2d2�E�΅��0+��.����j�������ܥ���v���q����X�����Ǜ|$qM- �'q܇�s�ta�u�'2p�Wz#7�Le��RUh���]Y)�(D��v���c[.aI��w���}f��`�7�z3p	����0�g�oD�&�0?��[J*BI
��IL�Tz5y�qC.s�颤�_�R�y��.��%��W�am�Gv��ҵ���~c��X�&G���+�{Q���c���ez8�ˎ�^[��+���1�!ɪ��h����Î� j�G�g��su�n74x���ޭ�!����l��/3fbǇ���J�tc�#-����t{ܟU�#���ٿ$e�\#���mk����rǙgEz��qD��;�OOBW�쭣7X+��dUg9��f&%�SX_�A�`���8 ;�)K���ȁ�<Wuou}O��H�z�.
5�a;o�̳�����BĦ5^S&K��nv$��h\��3�2.�NZ띒�("d��U�_/Y�����8ռ=���8�,�L�kE��&������N����t��kGG��P�W�D<o<��s�Vrk�[1^{���w~���>'�]����C�벨5�o#+��Sb�]�8�MCzl��	��i�V�k�����'+���K������9��3������WP|�&��/�땝gr]���`�[;�$;gfԸ�_���`�lR��=�FG����d�5�|9��֑ˇ� �ѹL�(�����#^k�߀�L��|$se"A0�$��=c\C~�uuą��1��ٙS�Z�/�M����rs"?�K�h���%��I��s�I�S�%��B��<j��N�AIV�E�[z�����Z�������"�;B�	dweq�|w�D��9پ�ЋYX��ż%]�۬x�y)���ꢤƷJL7w��`��{Į��`�� �,�+Y4��YY�gZ�@�T��Zaa!n��~��O����T-����|xX�7���=b�;�ڥ�h�`#�Z*�m��(��`�����N���17p�m!��Q)�q�g� R�㯏,£�ƀ�φ.�!8N0U��	���^(�m��\'�?�P���]c�h�����?\�|B����	g��ͭ�Ƨ��G��b�Ճ�y�Mw�O���y=��0"N�̫��Hk=�~]ҩ������I�;t,�cҫ�M���JiB&��H;�̕����`�a���"y�ƣg#g�k��1}�

�W�7�;ӎ��Y�͕�~0 �;��Yd��&⻯p�R��5�pq0Ѕ#^			��IW���L%��{E��z}B�.<B���cPd"C����������sq�@�9� �?T淰��b����Vt�+>K i��ȧT^���?�*+�/s�ژ��L�e)Yb9�苣�aH���ȣ��|��Pa��s��颣�J�;:v�$���t�DDg0���j;z�L�p͵��p��[���33��
@��Ą^��A�&u�������I�<ݻ����{x�g���I5�B��e��$��Ջ�<�Q���6]iR��`NH��$�J�x�����$����xjtַW��d����|���g��*ǂ4H�5E�Ip�k���ja+��&�k�G��W��`�¿�9��c�ůCD�_@��)�@���m�/ӟ�ݙA�VW�����>fD�����	<��.i퇹-ގ�P�`0X��Lq��K�g�?��R�Q��ǝK����lY�+�R{5v�aL���GHr^>7iP��L)Gb	 .�C�1��="]���:(涓o�>�I~GT���HҶb<�"J����o�:吨�����eP4$*��D��$8��R�<R@^iy�55t8��྅����$	ô7���Y���5�޼y��+nxb"�����p!΃323[��:�+�����M)�<�n�	��v\��R<���^��OK���h���j�:��Vt&��nI�b9���s�ŝ�נ�$�N�i�ެ�<��^����.�}�j:I˾^'N����z/�q0vM��y�(ztgG���$�3��n.;��2�~�vI3��	���C���ԗ%	�W����.�}o���#'�fz9�0Ш��-�ƥ��h[��;k�L���q(z2��8Z�����(u�!@ѵ�`�čj�ێ�6.?�50��b��,��uu�JD���<&��}�=��ZP���mm/z�i�����O�3N�H�`�L�݁�����	 4А���>�䥆�a�m9-P�M�+�oo�#���ԯ�)�m9b$Z��hgq���]�&)��܍g��y�O*���%s"�6�2u�a[ �a�.ۏ�e�Ɉ�������7!��s�Dh��N{��?1�[�YK��ޙ��$]dX'\�U��>�t����ר}���&tf�S�<�{�|Ձi4�L�����j9Qa�x���bp���YJ#��[�28;u��ݩ�� j����ׇ]��eŅoޜ�p͆m]c�N�'ai1I[ާRcK��� �^�����0V�L�{IZ>�q:jq]W�q�}�����N]��>�q�]
��fQ��M)ymM����.�CW��xYK�{k��^,��Y��K�}��`�����QʂH�D�����x�e	�����Prֻ�qI" S.)��>9.�Uۍe�����2�\��>p�P~\z?P4 ���t���� ��u#3�9��7�prb�G��AZ�_������H�?�?�4f��Ru�"��f��Y���￞���%$K/'���3�N3�/P�]�{�s���涤')�q��x	^��c����'}Ώ i�m�N.�,��@��A�Z�Ό35�m�[�]H�$G�r�X�0���TyE�����#1^��z$�~�ߣZT�٘�O�����G��ЯJ	0�@;�K��dK����#�&�Y�M�F��.j7n�_��P�PI�
O}{m��h<	�>�n<u����
zg�@C0}���Ks�(z����ZѪ�.&�߷�4�����3]��hd�h�k?��@�{_���ge���(�Q~��`�ԗ:s�e�C���@�
�6�_��J�i��񙮁4�������M�<�B��Q���#�p@�Їyܔ
 �Ē3Jb����H�ƞ%�5<<<��"���Pk��8J�^mRz��0"e?�J$ć��$�MEM��LD^��V�lv)�f3��V��fj�K�#p�����i}�jG��.��t�=
D�
���K���������)sF&��ϳh��^���~q�	���3����q�}�p�@[�UPPPf����\������D���o200�ʔ-3�"'�������P���p>�%M///�7TUU}��0j���e��N'|ϡ��d��¿�[�1}���@��v	����o2�=ԕ$g�ţ����gᄑ�R;���o^{�$�v%��T�DJ���6�}h8����:��7�<��؈�8�v Pꅖ�FP��钮*E>�:ύ��k��8���~��pV�Wӵ��ܱ��S�Ò��ܚ����S_�p�|[��2��/�Y����G��{���y2kx��xb����)���iӢ�������L��4�͑ۖ�7�~h�l�"�///ŝ�_d��>q�	��]����jҙ��j[Z�#X��-w�T�ۀ�&��s��"{�Do���m�Je����JU������օ|%��/r����WC^;�.�J K(��+���%����Jl��)1��������_q|zKy�Z��'nó�jl2w|w��<�,���-ǋ�b���&� �}�u��}y���c#���<��av������� �.v���ϴ�~�W~q0S>���=����k'c��߿_c�D��`Z<�Ԙ5�#q?��\snn�n`	s��n`svrx|���G�D"u��%lmm���ɳb
׃xĪ�	��u����(%��=�5�H�7U͒��˃�rv:����4Kpp(�$�����	��A�@3յ����O��@`ӕn� ��w;/�d�O�v��B�N���"�@��>~��bꍓ�#K���]K�=�w�b��}~V�ꥡ���^&4�pt�殕�nx�a��OW��:ʯ�:�$��2������i��g�d�,�>�e�b}���;���̶iY�J�^�-�
oy�!���e>�ܫ�v�9߳<��$�`k�V�?8�w��s�,���џ�'l�Q����?[���s�����{yM�	jW��d��R� �'���f�.����_��W���Z�5�\��OZ�����L�,�{�\�$y>0z��+x�ɪ���v��������`��`Y������S�5�ĚKK�(��R��{�G���3�v�:��`��7وSb��e!w�Z�V���O�{�lư[�沣���+d5��t�����/8H4v��T�E�	�+����/<rv騛D��mq����$8������ۑ􂝋�C33�11�m{��S���Z-�%j���⚛5�_�{xT���<�Y4ܫC�(P� YH6c��{�~k�.�����`#"���w�x�zw&�**�lS�o &�Iy�[�?���%{]u�r�j7j����q���-��y�񍏖�������%�&o16��Ck}@^�O;3���>��/@q�$	iA;�k����������4�ާ q��n3T¦��ۋ��$S��b�K����̪W�TGB�2�v,��oz��-�S�.=�?������H0j������O��Ĭ��s�]�㝹�o�W�n�R�؄� ǈ�zp� ���Q.����3��E����rvB��/-�����M��)©Ԇ����}r�>�'8��t%GI@�2ܒ�V��CR���ٷ��A�+�6�"�(1@|����|�����O��� q�ж���iFpI���0(�9=�?�  ���!�j�`�,R^4��``b��?Qe�^ڙ�}������]�
��(���744�y��TUW;��R%x�O������d���PܒK�^RcP?��6��h�Dk���Vdb~�q��է6��6a�h��K(dٲP�x��A?����r�OS���(]_޸8�����K��DoT����l�E*���gu>�7Rڝ!�b��X����~�䄿tO>X3=����f)��v��ɹA��˙��=�t�b�c���[�c��D��D}m��V ;�r����iX�e�g؍���##�DXn,9������D���c7ww�Ǝ��[�����C��(z����/Y{�8�=m7��f�%��wܧ�@OϚvy_,貾���릲�J�RZ�{��W�KE/�뿲����G�P<etv��$��fb�V1}(���m�R �:�L	kF9[ x5�b��psE��0��.�ʍ1�ض1Qx��!�w���܋�����q/�-1�c���9{�"��������2�&qO)f�=��S�\�<�"��m��	B�pw��XYYu�l�V���t��j$��)��cr��~Lf�s��-ҕ7����K3�Þi�!h��RE�Q��H��l7:��-���Zk
_�/�����>�Ը���A������y#���Y=�}���1��B$��鄹�L��lI �'#`�ORMԍ�
J�a�ʂ���vn��vJ�F���$��J�K��/3n��֦!��J�ɣA��$�~g��㿍@y��<��Q�7�p�5!RL��7��X�Tp�׫�|�Q�n`��ϧ�[����Ɲ��P�����v�8��W9�T(3-����m\0�OT$����r�����K.'��$?����%8�����/��Tˤ��R8�-�4�9&���o�6��A{�U�S}���T��W�0�2��N����r�O�s�_���P����^!G�?�݈�t��iQ��,�Ey�
jx0�2\i�"F!���l���/]��`��#&-��`ebaA����'��q�yW���qW,�Z�Y GFn�-��Fσ��!�`���ũ����vv|	�z55O_}n7�Y�5ITΘٹ��,�y���@�l;ۧ7�o�h��l�Ȓh9�啙k��څ�q����7�7m:#Ѻ���3��Aj�H�����uC�b!'Atx}xQ���؎�]΅��eex�MG���`�38]�iv#"u�~㾔�4_�m�X���w��[���3'V�u�O��D�3�eƿ�9$sM4kx2 4F�\�>"�pF9�x�������<j��[Y��<�Fb'��Y�4�P�#����{�cc: ��a�Y�ō@2�����w	���Qs��xx��)4��aܠP���`܍'��^-f)F�9-�YI��2 ���!�s����A��98&^�j�v�3��T,�\�vy�f�[��o@��_�y�$�(��з�]k�rB���G�g�dսl�z�an��;���x�4� Z��Ms��x*�V|�썄W�/�ˌ[�5���<�{��%j�fP�?MG�v���N�bbGǗ���^p������PiR�--�)�>LKKK��c���N����)�� j�����wB}q~I�K8\R��`���9d}=#n��ή���`hr�g;9cn`� ���pD�� ��)�J�,u������S�V�Y�VR(~gu'���W%���@K��$�y����M*�?W"�g�+�*�\"6^�Y��{.m���ʟ���fLN��b<*���o��d~M�3�p�9�����o�]��L��]p=|��K�ϴ*N�~϶�<Y���7~�$�:�~V�R?;?�j`Pbrx}!�E�&��oT��s�1���0������UT/��N�x������ַ����Xs''ʶ�6V֎�Aʐ��<EvI(555�G
4�������H���4�'aU
�RK �����ݖ���=�}�N4ų~��Na6�q#v1�v�[�zҜ�u�����S�')XR����z���r��3ukx8Ť�o(��Փ8Y#zH�ɝ��wz p.���[�1��B~+A���A�Y��3����zw㿽5H�,���������cL��fmW+�{VP�8Vvv�BQ=N5O���\��֖��߿I�ɭ��4�]]��{{�m����o��wW�_;N�7���������L��C��agg^O�<� �ITT��h[;;܏FGG�lRG�g6}e��I[t�=���S��u��|�� �A<|�4&`�nM~^>�Nà)�v�/j��04u��\:!�t����Wo�6���9����!xyZW@7���֍���b��RC�&ҹ�V4���3av�� ��s/��1~���Pwd"RT�_�u�Ay�q_���,Z�����rb�9�R����w~���n���X�	uf'��f��.��/��U�����l��{�����}a`g�g���5��͍&;;����p	?y��9a�|�㮤��p>|4!�XvNNμTMUUFv���������I�0k����W�2{Bb���5�C�w��\�C����Ip#�dP�)��������27��I���Q����i8a���%�,�Ʃ�dt���B��`|{o����ob9��>����Ǔj�I*��A�M�J��� ��Y��Z�}�j�2�_�6A�w�5/A�Z��.�`����������{��k� |��1�������T����x.�e���=3�}�n�ck������^����6�mn���S� ��/3\�q�>L[v�ل61���5��ÏO���y��B����&I4����o�����Mݐs�M�`�_�:�B��~����eT�;^�%W�}-x���0������L~�N���rCc���L���b�.Z���^��b��M?j�L}�M� }l�p����F	�c���)�|��H�Ph�8Qm���	��{��g�R���L7�O���̓;u�� ����[  �����(���v��	���\�4I����V��%t[�z�Rzy�൜��ȝp ���L}|� �V��)�231��T����K�|O��n����2X�gb�R�hV��*�1ڦЃ���TZ[k��ϖ�f���b].�Y��$���I�D���'�4%r��:OF�����GY�UR�����(7��#Z���xCf�[i2�D�^!Dhy]祊2�q�@R�0���ev��v�M��x�� "4ѧ_�wc߽�"XV��Q>�9؉Vg�Y��K�r��օȿ=�+䙠n��3���h�g z<"����-Ƈ��ڰ)�*�1b��{�6bNuk2h�ޥĜ��1�I.�.@�2[�/�17�eB���S"Ω�Z�n�;�H�آ+����W��X�U��eF����+.Z�*ff��6̍T�ۅ�$�)��cܑS{��r�i�;)��y�3�Ky����BwG�����#�i�2�Cp�i� ^�\oU�r�q(�K3E{�n�?�����"�G#s��.
�g��;�
�� S�h�mV��5�ev/v�)�eP����hR���ڃ��Q��-��gRN���G��M8��Y/qGrWGYڋ����Q���iVaֱ4����^C2ˎ��A�*��"�Ww�2��-up����,L�u0+!!x�z��B��-z�^o�*4�r�R'�9o����D�g�怯�*�}�i&��[�ۄ�\�o��������3�z	ѭ_U�M�Tl���Op��F��^Z�����LU�u�5\��_,H\,St\2�d��t8�Y!�<���3����/�������~<�?���D^�Er�d0�C�h���}��o86-_SJ(W3�0������z2�f�
�R�L��c�� KjJ�w�C�EWz^g��-K�t`k���X�N�����d G����}��"��ڦT ��?]��#�+s]��Ƥ8L��#6
��'��p{)�ݎ�j�v�]��b
3)�V�O6G���O��ud8�<���gb���fa)kM���R;�mq����-�Q8�Ӕc�>d���f��a�(�I�Zv�c�^�<`���큺�W��N�Y�2Vo#��V���뭊�3��
=	?�O����a���:ϢP��y�E�.Õ�8t�>�;��1�{�-k����-6�cAq����򞎕m�*����l��Z�Ɯf�Ŷ��!x݃G�UA(��;n�"AC�����Ût��u�"3%İ�����/�'+��j[^���&��%�]��4�����^Dl�r~Uo�r�-d��)Q�����bgI��I�1�چq�g�i/���E+nK��W_ �@ɢ�̴�z� Y�}��	��n(��=��E�%rn4L�������Փ��f�.�0�G_�8���?��O>}~1Fr9v���~��A<w#=�<�l̲�݂
�9�ŐQ�a	�tzAE�x�6G�u7L	�<��o�4N�z�9k�� �Bf+k� uիUk��z�Ս��瘸��׫eKH̦?��Y>�O��c�/BpGŠIak�w>)������8b��Χ�?��ç��� ���6	a��;4YZ���ְ�ٴ������}n��EpT��R����8(u�
���<���,��Z��`����Tʇ���9��nJ��I�C>��x.�{�*�,��8�W��X$��ίmV�#Pv��c�C��z\M�5�@f�{��\ʓdr.r?�%�U��#O�����-�6�OzRT]�&�-�i�+��O�(w���vA��z�K����[����碌��I�'�Y��Fr�-�W��[1ϳ�SM�GjȦ<��̈́s�A�"�l
4K�1���S�֒�fFj[�+l���I��R��Ty6���{e��|��3�e3��-��T%�������7<3��Ŗ&o�������>'2;���
ӱ��n#Kg*���3*�kv6��E�RyWy)G]�Rj6K�Fސxh?0���?{�JҰ%�`r|�2~�lNX��G�Z��$R�i���g��ih�0d�ȓ���IOy���0M�q�F�����eȆ\&� {ɗ�ٷ�j#��p6���0w�Mn�#�z�&!�:����,
�G�;�T��_� X��i�톇QϚ�.�@p� �8|���,�Z�v=���C�St]��. ݀]�|7F(�ܣ<�2�/ ���2���w���6�Q�܉{��Ơ��g�=ρe�<d�f�,�Na�.�\J\��4�s�|I&p2��]_EQC���1E�*�����]��EIt���I�QB���i�M�O#��eRj���}
s��>���Z;DJ���0K�(K�E�L��O���\��7�`��\��
I���8�E�=0��	G�w��|kQ����i�y���ʗ
h(��h��İ[�N�@�t	�/XH��.�����h��g�z�`��U��u�$��T�q��3BK��#g�I�`��ƩǂV�)�!q@��ئ���kN��=N�x}�sr)r��K+!���&[/�p�?��6�D�)с�,�M�f�͍U%�( �`�E���+:����`4���B���������%�zUʷW�i��in��D#)N��x�h#�uFk����x8��*ulIg���/�?���� _$�L���w�d�8����S��f&F>'�|>��ǃ;$���?��N&�
drS��~,�i�٩4j�i��o(�������	��*���/�FR����k��0��-Q\Z9+�2��q����!��3];ǵ���pD��U
�7��3�T���E�����X��|��V�W����3����{�H��-�+��tڑ�EfhB���1�D�eW�ƭ'e=gH�qI�?4���>}�}>�n�Uƛ�[�����e����]��/�M�~�����fu��׾h���Y�a���jՇ O��<f�<( X�`�zs��8N!D�,�]��>c���c�����#�b�I!�(��~�C��Q��������$<dUgV�|Wʓ�qH�%��u��GX���}�ϲP�Y�>Gꃝ8����g�4�z_L뼲H���^�x�7`V�o�*Q�!�ؘB/���8 -�nXq�Eg���c�ok/�nSu2ɸ���QC��Ee����&t�&���T%;���>8$�@gAV�=o�Gj��L��g4R*(���=���Q��k��s���u����+�<WǷ캢�袿u��:/��w�A�Ѿw&���s��nCL��޷��L�m���*��P�l�^�����(�)���%����ͬ��e9LT�4ʇpH�}x�'O�u}�e�I��S��Sy�HO��d ߬,���븡j)�}�-&�V7.(�'\�x�N�>٢{8t������k��u�>��X����La�y�RZ��TQ:�A����լ��b�l�r������Ѥҵ��I-���@���K� tAAE������'��M�@ �T��ؚt�R{�9Lk���U8�j��E6G�ף�S�Ҙsa|��C���D���P{��򩓬A�-g�-'���=u�a���}�%y�XϢC��,��s)	d&ݝ\fwYD��c�a2=��Œ#x��%�c<����g����no��ӮE����;ʻ�78���W �Y��a��}�yZ���.Y�^��7A�B�HٱST+�A�QT�1v��{��
��f_�t�Y�M�P�������.S��	yF��D�LH���޷C=��\��:��0M@�f�]ǌ�XD�p��O�@B�I7�r��<u$u��[ʾ���=�>�K���)'w<�#���6�^�cΟ��������Z��?	���F��
�&l�J�ަ��<o��i�aW�Y$�a�Iԍ�%���W[wI�;��j�D��e��V�o�o��C�7+��/��R=�~P)�����^�Za�{����KE�QY�~���l%R�P�H]X�W|�88 �4K�}{}JF�Pʭ�����p}��-6�pm�[s|�e��*j�4"��� �Ir��Ii���	9�)׈�y�M`B.��gq�z&�{����f�;uP�8�=-��"W%�}I��ӛ��s��p!�hST��5�M��Y�w�3�f9D�%�z���{<������'}Hf��|Bغ��=>��R�MN��ǡ�y2�#���+�A� k�	߄`T�)��ל�?���Gi��2\b�^��{l.�S�W{�y���ԑ�Ng��Tz+�,������ץ�Iн3/Rxޠ�q�A����=�����[֕%
|\��ꤝ&N�	7�ڦ�X2�u�o+��U�/�re5����n�i-���v=<�-��j@�Z��$�&�W�4B)�����MtȹG;�e�1���3Zyo��#��$�>�^���<v~pj�&�����_�f
�**�����6�ŭ�W��lF��^<�[z�~�xU��\�c�8=��hz������͒~�p�����&�����7�]�i��zA�l��7S�`g�U��k��,���J�Z��w�	�E[I�|M��[���S
�2WiWg�d5�Z��P���۪���[Sz*�U��l�Sޣ5�$����9P����+��,�2�}�;|���wb�AdIш��S,�m��w��N��-���\���ue<���+w�I�Q{Q�%+]W���A��Qe�w�}�@�8zv=�qjG}���w��V;j���(屖uQ)������������~�"s�ș1�6���"2�Q�{�z�$�[x�I���Gg�3�����+(�l�9i���'�s���xNɎ%�3 }��{�Ǘ�RҬ��5]W�����Yz��Ӽ�q9�=����^"JwE�-�(k�%M��#in��O��!q����q�G_��E7�CXJ��6�f��ϳ�F������vG�L�wţ��Wo�xwPՈu����G�6��p������;y�*��O׽
E!�y fl��و8cN��������N�F�����>}i�WR�JZ��@4��`��xp�C==�`u��g��E�U�Q��N�|�ƅ3ޫ�xl�+`c����x8S/�UEc��9.����� ��H�fg��L�z�!��bh.kBݡQ�/⎣{����;�L<Dm.\�X�XP�#KIZz&| ���9:c����A���&G훫�2^,+X��]f���E���ހξ�N��<Ҷ���^�
�����V_��%�<��^R� 5$�,�O&D>�m�st���Y�%�`t��W�S�P{�cC�|^�Ig���k���?8
���~z�`)���J��W��R ��^l�<����)�5c����M�;fN���/�ܧ"Dw[-�?r@/*|�It@�~G��T_��v�J�4�瞗3c|�1J4�NS�[N��W��hz���_jӱ�u?�rIe���^�6�k��o�9=��j�r�ķSK64ǉS�(P�cu�Q$Z�%ŽTmR鴢2f��K9��?�!��!A���|3Su�dō�w�7�~��oz+��~y�{H�t�<+��C�����-���q$k5�O������][ge���R�Bk|#����
�:IN�쭣��ma�{��!�~VN�Th�~%-0�ƹƴ^7/c��<o�`S+��L@��W�O�P����f1r@4jI��M��E�˸\���7F\��g�s�0%��!n�piK:!�@<�*W�:�2ڲV��Z�Dh�h�G��EhV�m险�?����%������7���CG�|
�j�A,�>���yp����S�p�����.���ڌ��Bi>��C,[����F\z�n$����
W�yD�bIhz�uӵ�ۼ��w{BA	��>׻��� s��5��c����O{��L��b�ڹ w�HRs뇹{�>��1�]'A̛��O��>��=2G]o��]naO��J�ٯ�[��&��pyd���) �.~���.����s��w�˺��e"u�7JRd���������t(;���%��zc��Vn�qd;���p}���$���#M���|)9D���|�u>ҋ���$�ն�)���<i�x�_��-/�R��Y������j�_��>�g�%�u츊a��V�uUg5�hSXDZ�"��̤�����xM@;®�d��\t=���VZ6���b��9��N��/��U/GІ���#W@~��U��z+�2Z���3c��w����`�X�@q?)Y�9%*{�hY��v��+q��>��o�3�ܢR����FW��b�!#�.���꥛�*�>G+�n�~���zf����S"�Ց��ZӛnMu�2�K{���d������0��eS�JOQ��U��e����JG�|B��d�����8�ki#�V��P��/�b�y'�HX
�vq�����������?4�W87�Aj{��'��d�w��ô�;!E'���i�)nЧ�x����m��I��%��s�NR�JV5��!�����ԙ�U3�ɹ[����[�XK��I�h}�@����%��}�6�sz�_�Lc����O;�-�(�.X;�8����9x�z9�ؚ,�2�ݿ�(��ޓ�B������4����P!oE�9�\ٰ��ii�d�������!x����Y�h5C	$b���Ч���8�&��b�p�4/�h/\҃VumNR��IU�K�\.m%�V�����1'��D��I#췜qW�ʵ�j5��/�w��'0k5��E��8zd�Oa��x� ۍg?�yI�"y�u�,���O~VV����`R�,��l��f�f�mo@���"�����l�p���_�|D�[R�4�ɨ��� |Ơ[% ��C�>GP�@=ݖ4�}�n�U_Hq���,��/�e.t�������:D�����d�$�Ąe�q�������[\����}�����k���2Jo�Df�J�ٯ���u\�=�<�����:��:n]�.88ː�8%��M�1�p��(��ϊ�Ua����=ü>����l�J4�i�7�&}�>h2}/����� ����fbd�e���ܡ��r�MHV�[>����[X'D��%��^�e���{��.U�>e��?Dy�p"�2
�B��� d�Fz,���.�TY�<ϸ;�DC���GW_J�čc�>H�Y$�$с�r
{���*P�QA�p���3���L���)����#���g�S,�y�4L�H��&7lO��HV�ũ*q����� �*&6"��$C_��R#�=nHY�}%����uB8�v� �@u������?�tB����ѺAs��f�+��^�HWj�3֏}�r�Q�E+�Dt�p8.s��q�@�c����8���x4�4qwZZ�K������)O�u~��)uL���F������� �]ze�K6���?����lw���e`�V����Њі��t�F�iq�"�_h+����:&��/��j�`ῐ����?I�P)�Պ0^�Rv�� n3X�r��o�ny�!&z��|����M�*�|��m��V�[�q#��|� 1��#���Xc���ms!��h�<>�* �:C^�)S����x7x����/t�KA!��	�(.6���i���ރF�9���ϳ�O���gL7��}�"u�'�[Ѝ�Lb�E�[�k64��?���O�j#����roX��$��o�M�㱯�w��r�H���T%p}bD�VO een������O/Y&�nr��?뎸�D��΅0�{�o�㰬_	U�Ǖ�p�ӄ�R����w�{A�ܶ��)E���jE��j�����x�ӒR�K��6��3p��*��̫�e:��\�[��3��T�bz����[�%����C|íO
�Qϐ�����b0����\2���(Y���<#>�V�8Y$��X��E����N�`�� fy�4u�x�<*��y� �!H�2�ϧ�'�W�����C�N]v)DԮg�ٙ�ѧrSN�QlfI\�"Hy�<�|��G�;����	����ra�-\�����J�S�Zw��;���-��m,xZt�`�3�ɴcJ��]��5lF=(������ʧT�R��������;�ex�
�"GO�Ai֬^�R����R���	�90�и����4���Ad#�P�Km�~ �JfXF��!)(<Uhg��P�L�ڍ�Q�kWŇ���[���N.�v3��\`.Ckn��R�������5C
>߹:0��wT����ϻ�0@�q5���~w���0O�d5��埅��ֺ%���9_���{@8g-O,1nS>sR�>��Ѕ�Ee �P���23}�:�|)��1�нO��h��Y�m}�I�l�`��
��E�Te��~�g�W����ꭣ���7P�iAT�Ni�����n$�A����CAJi�a�B������]��yך�X�����~�}�9�,_|�;vȔ]�ؽ��G�&�t�v��f�V���3^�����v,�r�xo=�-�i��һ��n?���B���B�H����@;�ү.�T�>�O��Ɇ�9�n�K�2f�$W+�*�>�	�fQ\=��R'�(�M�\I��η���v�h�<��Ag0+Zs֔hCXw�1b�?�@n�{�vv� <�y<i��ѺN�"+�!v��r�!���lk�p@��7�Q���E�k�=��ƿ��L@�H3ߌМO��FwH���^R��CN�#nn"�%wt�=����o@�-����}�k[�o5>�<���?|^^��H|��ap+�!K��2m҆�y�d�~M�Ē��+Ih�.d&��<��7���+�c�b���?G��]�
.���:��u�3�s�K3��q�dd$4]I���ϋo^=듹��}Hf�Y���?���H_ϗI"j�����`@Tc��񈅘3�M$�m�1��=���! �a@�u	f{��G�]�
R���}96���i���sQ B(���\�߈�LC��w0�7�u
 i�V��\�+�8mw:���揣�|�Ԟ��bXh!���k�=V�O�9���V��k�v�e����-�I���(Y��>6���,A���F^�����C��!���R�����'���'#�W�"+�ْ���b\�}$��d������VH���~S�b����iFş�4�h��Ӗd٣�69���.�gu��Z��D�ц��,�=�jrw��.��]cL��u4eY.�[�D4���K�+8`��wI����4ŉ�Y^�.�s���$
�K��o��}û�=?	a����50����"�
���$�!�����f��K�l�?�IВMm��F
��?���4�t��Z�-�d��.lP��{�ȖT4dg��{y�3������v�����o����R`�L&�˗R����/u$fj��-����Jɯ[�u�7�i� ����g��͡7Gh��.l��A�������߲�����Y#���S����(�����`d�-[�j�Nڑ�t'.��Vҹ������)qj�����pw1+�3���z�	΅��Byl��~���3\%qEw}��G���(���,Um-r>��BH��P&d�2����@�����8]��J����S���lw�/ڎ��H`�˳�^F���׆����������}�7j.�R�H���a����L	�vr�k��Jf��EJ�̱LŲMN�rjcz���)���. [��d���^R�K5�6ms��W�Mڴ����D��~�jmB7��(kBA��?�K`��a3�o� ��bC�L;���ܒ`�t��E����0�]D�n��}�{4� 7�#�a��ɩ%�T�!��!5�Pk�1"���)h����C�pZ^�Ʌ��p���d�OV'n��5ǋ�xOM^秵&��&���u�����X@�u�sg�>M�A`u������&�X]7�������I��r��U(�y����8-9�Qf�4<��-4�V�=��L)�%�]�xQw�H���i>�I��y�Ö%�$�W�u� ����`���
�����8y�{Q���҃U��<�̘;��sꁟG�tZѿ�����O��;6�0ި� !�;�wH�<�m4��.֬��nˣכ2~Jg`Y��@�ö
Kx���ϕ@�W:-�9U�{�1���_V�:��^КA?�j�=��$�/�1n��K��3oAZ*�QX�\�������/���J�����}��t
p*O�&�ҩ'���!0���H�ےc+8�NI�����;V�ms(F�S�r�R
h�m�zR�!H���~��ZJO���>�� �ݺ��Gǵ"��lgK�H~(������(���x�Gw��A����!�1J�sD��3j��IҬ߬�Q���U���r8O��z�^�{XR���Z���Zh��0��{�#�e����P�6o'	}�;�`/��j�yL�I	Y]�Ә�h0z�)�I�E�������x䤪�E�c�14!ݣ���n�p���(qU��9�56�t����"� A�w�������}iԢ-e�-���?2F����!^ǟ,�4U��j�l�M����^�S���V&:�V�D�����a����5H��~��v�H�LG,��>$?��,5e'�t2�N�/�m��@[����:��lk\lc�d�-��N�^����� [�<��Tv�w�g����Q��$�?�i��'J�0|����P&E������j.Y6��J�����^�J��Si�2���+� Ф�'��D|��ܹ��z���úN_ƛz���j�>A6x?��8��nxӺ���vH]� �Zv{����/�&�b���a���D-�3]#���xa��x(�3�X3`��Y����n(�$]8��;!Oֻk&G�)?yx�c=܎���?�C���wY������ag#�,��xz�M��&�QW?��%��6�J�]���w�\��(��`zu���{��y������Z�8�c����-R�Ӕ���ݔ��z����:�F�!g��!D`��&�!�(Ύ�F�#u|�; ��	�/VT	N�g��4&����Q��(ѕx�'2�3z�#ch�Q�䵼��J{
���w�mA Lg���I����J#��L�c�o���#�׾,k�Y�źq�{2�Ɂ�����z���>e��</ol�{� ��eq�t�|<��Un���T�Πz�*�ek�4��roa�mj9�\p�c]����2�W5Y�m���Dw�d���$|9g��]���/w��>�?�Ń�	]�V}�+�D���Ÿa���6���:�1Hl��'�h��@��3]c/eY�_���5��k���V$�(lA]��O/1-�����-�����b �<�����3��X5�:�:k�3ep�%5���}�ɿCn�S�;&9�ߡ��2�O��oi�6�����t����Gfp��.�[�gAa��s��������"o���_���F�<�>�gU�J�v"j����
,��d�*�R8=��k�6����g
N�^|���[�5&i�b=���z=���ƣ����X�$�	���_��Ҟ��I�~b�W�{p5�lK�ys"aruP�!?����l7&)6Ң����)"�=�7��47�~����\�����"��ގm����ZC7�ϖ�׿Nc�3�!7ߙ��e���9%U^_��ɊȄ�<ޔP�+�֟�o��S�g%I������3Z���GT(~�I}��?N�ؕ�R�?̚��栫ߨfwJ���Nt-����{�J{E1PCot&^���$��o�b1Y�n1������wx����==��X^��7O
«��9�b��6��V��}�n[z>Ps�`�Փ��l2P��J��
�J{n��@��q���ܛ�F��F�P��H���
~ .,�)�s���j1��n3�d�J1˖�*�匏m2�;b�f��V󟗺����h�������ˮ��
@�3���Y�dJ�$����t#DD��OmO�b��X�j��~�r.o#*�	giz7D\ra�������:�����������Z�F:U��ʊ���M�|�Ws���:�!w.g�Z�ۺ�
�1�)Sx���a��?h5F^ D���7�X]P��#)h������i�1^I0�$$4�dY��k�vp�>�Y�FLy��] j���W���>��=)y�q~GSL'�Gmqvt�st��"�C�����C���`	?�i6,�I��󛲪���A)C�I�>�
����eFW���i/̜=,�)�����fݬ��쾮�fP��F��b��#�^X��;=�M\������`2x�[�$���4�{#5A����������2�.I����2U=5�Ͽ����e�:� Q�ok'm=��n�_Z���pj�1 a�:U%}�Щ*�I��5�~UvD�5��|�'��G�
���OLrf���=�.����ZJP#X���b��Zyu ������{z��>	ʃ��ոG?L�G-Z�H)��i����AS�Ύ�d��C�G��dU�}�1B�|<��	N�+X#�&㉤��}K�� �\گ�_2��w��]~v��3��q��ӳ'k��yT�'[W[O�:r}7�� e�u�2y��/�.�l
@������.a}�]���Ao���n�4d�S;��*�4̝���>@pN���y`	���5r�O*����t�{y� hI��?i����$���D����n\`��=�2+��/g�^��n\aoi;~�_��Fd��^�	�G���ꄰ�p��Ə1ׁ����9r&��̺_1 Cﲢ��
&v�L(	@L.���%W�13���w>ZO���9��(DK���"7&�i@���ܿNys�fj�w ��(��g�rnd�R����8��:��������>�J ��Zh���h�Di��ӊ=T�7J�{��.�(jV�K$��!���`��������3"�.o�"~����ڤI���vlN���|�0Gz���R��:���w��00���@'�,���!g��ى�-�TI?�l�����s���O��0�:�F�����Ze���_+�q�K���WM,ڮ\�5�ׁ0:yå0���Vͳ�%��Gã��$qJ��x��]?��I� �^�_�+pt
!d�ͱH<����	�W{�3iRS�/uq���F��u���%��(SNJ
gB��-N���y+�}f}�zM�Pm�6S��n( �Ϣ���+�i*��g7�� U��d��(���/�=5� �WJ���kp5����K,I�+�׈s=?]�Ճ�z�q��qbF?���;��3)YpEk�p3B��ތMR{�:��d3�x�,?�����s�@���Z�aw�mwh=ȡ���!���V)���`Zntt-��Ώ5�fw>������o���4lm..6bBjQ��ܔa�9rt@�x�d��ۋ[wlOY3�l���5���7�
���h�Ǉ7�p�������r��?͹O]H8VO���vb����W-��L:�*�oT���0�,��W��ߘE,{5FF����<e#j���P��>�5.U-�������g����1���@�{ZMp���f\��d4٧���y>�J1/I_P�D�1z�����m�~j�H"N3�q�t>Q��ѕ��5b,Dkʄxy�ɓ���똌�#�ǡ���t��"�(�~տ:mxE�MH7��=����Qt��ѝ=͆2nD��QKɆ=�1�UKör�'��qJ���
8�Si����*t$o�s��:�~�֥N�S��4d�p�xD�A�|�}�W����W������':�E���FA	��o݅v����{~�K���z��#�(]�J��x�t��	e�P��~�B��BP��Y�9Hj7V��x6*g'���\����>�U�}��5����_���<v��סZs�ڂ�T)+L�AM�~PH��/�����u։�j��y�?��Pb�=0 �L ��G���k�������TsR�t�p��X0a'�}��4I��T�|ND<i�7��Fo��������|7�S�y��?)�$�mk��R�L��Z��)���z/S�o����8'X��G�6'�SQ2Ň�iy�ks�S��&���Ƌ�߈|�v�3��{p�x2�,Z�/s�8����b�Z�9!��\N��������:{�s���~��⹘6���2��&N�{T�Ē	��hV"�W�}���r�HV9Z�$�*��yֿ���� �Q�j��I{���z\��%H�Wx-�7�wLKV���4��8bQ�j�L�<J1rq�o��<�d�\_¥������i@�����#2���"��Jj���]a�%���ցB�Bȍ��K�E�%�/3�a��E���뎌�ж�ݻ/G�m.�yA����?� щFD%�]Z"�mda���P���"*$`<�� �;�9m|In;�1�{�5�&F�Ys�M[8��x¸���ސ�1��}z���s2ȶ)jcfQ:"�=�]~[��!��];���d������?��l��.�����*���H����a�����ݸ"����<�,��s��V�\���oO(�=¹��,)��J} q�2o�����>9�)�|BA^����cjW�xC(�æNAa_���md �_ZS�����|�j���d�|�(�=��6M��!_W�o��ۜ�a��@՞�׋�෠�bv�`�Q��_--#K���9\dt�j/U;j�Z3F���]�����o_E���A[�FQz=�&��[r.7�9�\kG
�A������:X�`��~����8�g� J qx���X�J�nb�_*0aU�m��3?_I����,s�I5ͼV�z;����^��3)�x��s�V��K� �Z��?I���.!b;���+�k�R"�w�jċ����	��I'L�)5ZT�0�F��=�Fy�����o'���������� �(SB���D�##�;T}��v~���P���̹��/�������U���&�J�^�ނ��?� �.q�Ʈ���>�)G[�ϻ����LGke���q����\�ӍSϔ#X�1�U�Xr�1�Fɱ�:`\nx_Va�b�̇��􊻲~��i�����!��(%>���o3#X��ʙ)���jז�����߄�[�wtg9U�}����.w'ؘ]����27w��(5�w�缀_7�U��O���h��a��m#���ϕ��̖qjG@��a�,����#���>���A�v�BO@L�dV�sl��º��q!��z�wI}����3l#$G,�8�{,�����o@8c3��A�?�����[�[�m�_n\�oJ�7�S�>��[�N=�!氏��iq��Z�%a�Vh�����&d�^�P�[��HF�%�f�cV��2��E�N���c��V6p/������l�a���[�/��a����������[	2�ka��k��f��;�j<s�E�}G�k�"sj�C��#��q�L7Ă���Ѱ���o��� ~QdC;L��w�f󏆍@ ���1r?r:AH�rCa�C;8�%�'�h�L�L����{*��o�@Dt�Ies���l�:�}�9�"�$h��t�NwRXZI���$�cv��ч����I�5͍��s9�B�~��m������O���I�Z&ݢ��v�U�Շm���[A	�0ha�8@���t��r�4�!6)g�L���bNyA�֝�/�s��^��ү|O�� ��L��*=�4t|��j* ���RxN*uŒ���}Q���봞*� ���v���mZ����v��ݦrM���U��f�1�����X'}��V��Eh��8Z��d��Q�Cf !���G�4��߷�`� ��R�{R=�FVv~7����|0Y��gEU���H$"ǡd�,��Cק(�74�b�듇+���>&7�IZ�MvZ��ڣ����������!�F�I'm�2Sﻡ��&�w�g�kL�I�����%X���װ �h~d�s�����H�מO�7*�a�?���YV�rw��8�����7i�s6�E �j��4���8fh)��Οz��׳s�p[����\�u�Pa;-���X	ZX�6	<�*C����H���U�	����-a+�A��H�@ta�E�n�ud ��z�=D]+�u���^<b�%��n�
\t�_ܛ�@�f����:���O�[9������-�m���su�B�TO .E:)�OIP+�G$S�����`/m-�I�r��'v͈��ڍ��� ��D]�Y�D� �Z�v��_P݀Y�cCr��g_�&�#L�8��'�>��A��oL?"gE�ť6q�N���9C����e�����ц?)���.���S�"��96f���;[vA�/�IF�����D8e-w��9���:����O~��ۋRL~g#��XO
0���i�y�RW��	�hV�ӭ
�:���{���}L����`��4�HI-ڭ�1[��օT�l�J�#�2�X�v�#��z���`B�6����D-���!Hi��ɧo�f1_r`�����U@j&M�YZ�nٳ
�'�3#
[���p��8E��bT�o��f��ƌJ����c}��O�Z�b�T��HK��E�8�N��ZA�&cu 2 ���FL6v)_GF$-�� ~D�8߿��~j���Ů>d�9����⮡8S<��3w�~=SK�	�.���Oe���X����oĽAb	H��x�J��;�N������)�ݢL��u�_d_�*x�(ĝ~�f���J�Ƚj^�N�,��Ci�o����S�#�f9UX�e<2�����`�طIe��.���x�x�<��L�iz��;�C7�g�ZN�Yo�0J�Ț�P���*Y���I�>:���ju���M����t�������|��)&�w:L1{.?����׃���J���S�_�j���il��c,�I)	��Ӝ@n'?Q�6��(�N�g��ACw�M�ly?�3wûQ�fT\�����h��T��O"y]�"��⫷�=�m�I��`�1e��m�oh�7�W��*�`���a�?��>��{Ya�6x�msSz̵V$�'�u?�;����w(�
(�hν�[s鶒D0pk>�2�j�[13�E�%1�qN�zU��Z5����U �)�Jg�K̳@�An��`�ޖ�:p~eX_Y�Q5��_�y���>kEn���&n!\�]��l���G�xU$��3*	����5��!��~U����q],B��n�釘�4�n����Jy�ދ�W��i�i�{%���J�[�,)0���Vꨇ��8�bi��8�JZj�O��&:��z��;��Y�)=΢�z8�\��f7��������\���'��I}�'�Ļ1����P`�7QL%v_�@{��{� -`N�G�0���}rϽ^4���q^9%M��]�q��ܓ�XHmPI����[�(�[�L�<���^�䮊ܓK�)�<�]-K]�߻Or%D1�')����:����;\�4���eS����`f/Zvx�B��N�����1!��B�5>���_�y��o~�\����^�.�SQ�JFT�M�#Cd�6����I�T���%N{S�A�4��C��rX+"@M���q�{'s�Dw_,n*`�?��-X���8�ͻ0�e��ۈ�ܖŉS��Kqq�8�j��l���
�à<�F�ԙ���pE�NP��I\�Waקt]��4��+��R��I4�勆.�����hN�8�~����Ĺ��I�4l���x���Z|��/��@#�W�q+�&U+t\�Y���� n�K5��jՐ�6gS��0�N�]"Џ�hգ��!vU;����i�*�0�9�c-�	��\�S�W��%�p�?�z,�8��Ҭ����W+���P<I��ȕ 4�,d�_�5 k��-Ε�i�@0��	"�OT�*[Si䜁G���j�	���%�AE-��Em���E��"O?hB��Q�.�虜v�` h�)~�ôፂ+�#
T�h�`eڭ��CV�h��C��,��,�����׬R���7d��%��?��q-�>�u����$��<)��G�;�8���H:�c/>,�+�減F�KUf�D�3�\q�_5�p,��/̕KL��zQ":�$�9�
ޖ��v��� ��tP��Pc���6	 ��>�k��C��2nj���N��T���B�=R,ع��r�*mRyk���q������¡�~�D�pt������c��f�k�Ϙr�/f�ݼ1qiH���6Y�sR��p�Y��R��i�k�[�֦��x)jS���"��A��DD�*�F(&ob\mW��ơ��e�3��"GkM�m�ŸMc���ڎA�Xn�˜�b�T����I��CF$$��9�q=O;�ݘ�I�4q�\����*�7v�Lb����)�N㵅$o ����� �NU�'��D���3Ȇf%
��Z4<��FȣL�n�R�J�mG��O�:��h]�5�y����ۦ�Ӡ�����^j?R9��ۍ@Gɦ�U[N@��Z��W��P\qY����O)~�FnJS��R��P��^�LƄBC�l��GSN��9b�(��=t��DJ$\7ǥ��y�����7���Uva0�vc��Ѻ�W�ō|���@2���Xe�h2�:ǄBbd��%ic�tZWZ��J
���ƛ�~mM)K^<��_N�jζ�_gn?y�,�$�.��dW/^�1�݉ީB��l�;���k�`٪
+���>9����O"�G�0&�5I���Gm�t4���l��"��v4��_����'T8���":�v�C��O�B�R���L6o�c��r�z�ދ��S,��'�}Wҏ'��Q�g��{I���b��t �k|�u�AS��|�_݆��_��6x�g���$����[_�kG[���i��Gw�1��\��J��K�<��*�S������R�N����z�Q��)LE���(T��~�$����G�
K�lN8����=_���|�"���ϬW���9E���2���|4Ԭ�9��ؙ~�OK�*K��F�B�D�("���T�iI#��?U�	�ԛ��w���̽]_��t`�x��^c`I�g��IK)E�L���
qA�)���]��\-�ϕ��g�Z։�\r�PM��Y7�Y�C,B���� 9	:�dϦ����9b��z��D��B2�_ўK�ܥ���D��	9�]��|h`/�}�{����T�={�9-<���%����X̽��1����|�ʅ���y޽ir�.� �цh�=�+�ɲ��^%@E���r���a�zs�wT�����͖f�;����}��c���XFt(F;p�$'`������Q���Nbt��#���Z��ױ�􎀝�\��Tk���}��'U�c	:G0W1��Z��W_ �QCU���S��E��o�#*Tæ��9�ϫv���R�ߛ�?�.����
Xǒ����-N�Q����P����\�	�r�`H�:T�v��R��'%F�iX��⽿����0}�ӗkH�#�$����4��?����͉�CF��;F];�~'��_�Zo)NG��i4]��]�ݿK��T����c� )E@��Dc�o��-�,ؕOIH" �~�;���� �7��v����h�{H?|�������6	�6�6cR$���*6D­H�ѐnŒnoBf+�2���'�&�s:Უ�%/v�}k��?�d�n�AD�O�n��̻	W:,���kY�>��k��Щʕ"�Nt�Mf���t�,�B�����0�_��k����%Xw=�o
��ί�:F�iHhTjIY�j�P�V��D�7�����}��i7��$	��A����Q}:�ɘ�Ǆ~)��dDkv�0a�?VĨ��"c
�;Q����֍��hːq��"q�:�f������m�]��(�븤�F���u��e|zx����Ӑ��;8��7�i~#Ɇ`��A��E���*Ro"���2]l�6�u��q��L�_`Σ��>��*n/,}���(Esp���w篾Ҧ�������)08�ײ������[o�b8�4^Z,�a��lP��	 ��\"�×�ĥM�hZm����,A۰mT�����4�`���E)�q�!Nr��F��0;�ٿ~}0p�8��?M�\\��X�DW��>����W�JN��*CQ��w���&k��u�`�B�L�{�����Z5���k��R��%�ũka�(�@p��A8^�%f���B�G�Q�����9��-i������>!7%j{AG�S1B�b���&��� ���|�<�]&+�7����}EF��GI�G�z�M�����V'dj�Xi�,�C�޵�˿��ތ�;߻��z	B9d:�Z!G�/��]-�\��&�xZ��F�a�H�_m2'81x��
���V�חJmp��5lI��T��\>�R}��9�c���YF���K%o��}��f)sR�u,ϒ�I9��O������ �2�8w�ܺ���~�v�`N�x�̩��^��Ǜ��|��7U��c{���O��4(-M����t����!�Q��,ȓlɞ6��qTe2Sbo65d��xC��Z�˱]K�+x��P�m�"�zF�����B+��[��k��
W�SBc��*�"�9M(M��X,#F�n *%5J� �Z :�}��7���B�UȲ�*X2%β]��b�� h���<����]3�@{˦��G��<U�&�h���p
�9c�{ڔ_����2�l6�%\EQ��3�D�J��G!����S��b��D�/ �7��3~���o��ܒ~��Ö�W�f���Ty�1� �0��B�9��R�ϔn� �sY�r�mB����gՐ ;�㍖�ΎJ����Ű���p��3��oķ��l��שk�m�J����Gof��y�l�a��מ��톖 Ŀ������g����ҷQ��&�����-�귋��+Q�gD@j`������M��<U���S+������Fj[{���G�5�o�%��ۿK�*C�$�)�Y��#V'F��A�Y ���F�%|����47)rq����j�E�\<�@V����Uh�ށ��V��Q��O��V�]��ɵ~��ܤ��3"t	��٠>׹.�qJL������|�}-����a^5��M꡵�����Ӣ��u���� /�t��'߆���Vd�zX�Aa���B����(v��=�tkuق���?�p�;���imWN�y�4(,\j�'���f�f����c�L�ɂ7�
^X�^�4�`�Avp��DF����헁���7�� ���1�>(\�ݹa�r=q���v ~3��w�&��R?K��8m\���V~c���z?��s��='
��M�_�6�;��R=��l���Oq�;�eͿߕҠ��	08��q	aR2��e�f���G�"Z�ӂ=���yfO�����%��)Ac������ʮ�������, ��9�r��I %ՠ&�O�3���Ј��'"�hco��i\�4��G�z�ZN�ݯ'(���;^�1|+�`���%����b!��Fj�SL�;���*����	�����7SNI�G�]�����bLm�IԖ<��S�S��J�ޑ����ם���mf�2�eCGA5}����g�Tk��ױ���ۻL(��*����[t[-좬�R3�:HCE8�[k��"T��2r��u{��ć��)��q�3���B]�s[����x��-���M�o�p�HH�n�o�s��ki]���՝:�x����U�谥z���%�K1o|�u}@��t��/��-�,5�A�Gѧۖ4�C����
tW�N��9�јA fo��C����:rqkNe�g���o^(1���D�cˤ�W�;�.gJ�"c�q�G�h(\n�B�Vo�.Jپ��G�]kCv�B�Ă�H�'!pGJ��d�����z\�QpK��JНᤙ��Jug�:������c�XI�UӰ	�[���e,0��!<45 �Nq���1����,����6� �"�J��V�IX��Q���)�G�ֶzz|��*:�� �aɀ�:���p/�'�I��j�$���t6U"����p"�G=cl3��܏�>\�!�n��w�o&=#ylG�n���Xw�%@(�PX�K�d_S��7ίv2ʿ���%�Hq� ���s�zɿ���9o��_�#%z\%I>W��ZF(����j�=m�K9+bM�F���,�}WhƎ(W��% x�Y��0�)���$�z����_�-��_������c�w��l-�Id���zp�n�'��k `��x�@�ߘ0��(B~i��(�j��WȔkN�4��"`ɢ!B� $i��Ì;@�����!\�|g���b��U��.O��u��+���N�Ԡ���|�u
�y���M4>M�ʆ�d�v�~�G���`h��H��p<�t?�	J�N,Bz=6��W��TqH�`~|��@�FWa�w�OS�D�	��4�4f0i�-+�f�\���RӲ])Q+�k�`�+	��>7��Z��X}�i1���˧�DbS�ʛ���_��W�(N�S�߱���%-�Q�d�ŪW�:�Zhg	������7֟��@�
�Yp~�DЕjP�׬XZ��>�z�f�zW��E`��Ί���y�����::t���p0Ư=DpH���%:��}�s���9Avh���L�a+��ٮ6n7WC� 3%��~E.�t2��\��2�� ׺G�ّA��4�����.�c�g������n!���]3N-�<W�~~&(����p��2(�0�գ~;خ5Y*�j7�ok0�6�����$�XJ� 2�y�Ibj�n�H�r�N	aO!���QV���=�Hr�t^�Qu�:�M���ӧ$�HZ��{N�]n�x	��"^xC�|��+��O�z]\}�	����?��OS`d�x:?�����d7Ͳ�,��]97E��n���C��C��:wcF9�u�hi��z؋*YK:hi1f%��ز�-��R��h*{iW"A{n��豚����xo���sRSק���5���rI��H�
�ƕ�[�zu]�W�c�\�J�/B��%�q��[�B�̗��z�X,,͛�*����ii�8����Ģ^��j�q��B.�`�1��!�۴%RT��Ê��2 ��~��KC�#��\��I<����Y���E?y��[	uX�T�.�?�3�Q����Ǆ����q9I%��5�f^�όS���M��DQ�]_T�iS��P�̷��j���WsM�5
��4�u��8󇘽�]����*iC�.��=��k.ب���Iy���:�ߠ��ݡQ�y���c���%
O5b�\�׀��/�jۍ�%�y�ߩ�a��i���S�]���Q�<@b�LC���x��I9��|�:�a~ʰ��;u�s����R`]^���PSJ�x@�������m��s�O$
+8��A��4�`��@���ʙ��ظK�s�5�Rn$�n����h~�kdУ����{��~�!3%�2!�o&��FV_ns Z������!���c����'M���� �Oh�~n,�a;_g�Z��r��Gp��oA��%#��� �~��Z����&K�;��֮쵑 S��]�y�uc��i�ӈ|�;m����j*T�z�U�2���<-H����im	1�:�g�"1Yr)Ӏ��1�-2�_)� �-E�U!O7zY.^w�/)K<����Y�]ٌ.M�F.� v��u�ѓ�[7�]�3��kɓ��u�+
c���/kq6��
����Z��;-%@�.��	Q�ֹ۠W_�!Zd�l?F;i�ƹy�U���Nb���2�_+7��}g�fp�����+p���){�f��:�Z���eX�]��|!7�(�����+�+lC�&5�y�Y0|G�X)v���v �]N��៱�(����~ƃ�Qf�A���2��)A��,��Ja��^��7i��	�)-�?9`v��'�7띾���RŊ���c�����Ԑ��}@������pj�����{x1�Y0�D1�y��):ç��d��q_Dfh�d+�^Yh�/g��A�u!2�r�M��y�V#���>�0��m����ѽ����-&�u���*��x��I�jB(Xܚ����n;dQp��sH�&����#(U��v\�4	���m���1~0��v��hw��XhN��ş��"/�_r��u/�Ē�3��b��EgM�a��dM�2,���i��X�G^B���ޝ0!Ԏ�Gz~�z�'�M�Q�D�}2�J�#FUf�80��?�xa$�~�~V).@ ��dJ����<ٶ�L�������h�{]������s��R7��쭃��pU>�ĭ�>b��1pT#^Z�EYZ9�O��y��>�{r��<s)A�q�%/M�X?B��!��3>�&�Ls���h�?�H�Cؽ���%��e_��-��!����A�7� 3�-�]Hoo���BkQ�1���S_=�(�5���g��K�2�K��ՂQ�x\��.f>��+m����wG,�/���Ŕ7_V��31�3�Ũ�*��W�5l�{�N����b����i���H%���j�e%>zز+|�f"��w��r)T��p��'2%h�74(f�_��n����J�ѕٞ<{��"��I�f���E.��fp���g������t�^J����6�a+{t|�8h_[��S.}�����7EKV�p��絯N!,Ӻ�wñ�ݕ�U�˪��3�����}��O�^��@�*L?�~�j7�����(�:���%�Y�L|vf�F.����Q�eƪ?�=+����TP�`S�\=�P���J|'��mN� ��[A.A�X�(����;��[<X������x�\���*Au��"� 4�~�16	yE�#'��:�7#�O�C��W?x����<+��f;�����S�jif�/�
��S�z	׸8ÿ�֏d�c"hɞ�ڢ��+
.��.~��NR7�z���Z�}8%bɸ����u�s��(��Ά����ej��t��/ ��ҫ��2^�(�b��^�q-�tc�P�!:O��r�@�zG��ؙ��3�~䃒zp��:&)@�[��:�LS����{����TȇEe,�Ą�w��)}������/��͟~���������}�:S��J}���$*��F�J��?d�T�]�-LKq���S�]
�P�ݡ8���-�Z�]����Z܃��~���ެ�E��9{�����<	���`� u]v5Jh���m���"Y�Y�ra��(:��d�$Ƚ	�5�7�D��M/6�x���2@���zcj���K����G)�/Ǎ�*y��#.rȲ~��S�;ώ�9��ʼ���K��@1.sD���3-(��o��`c�DА{�?d��ۯ��	"��6��-�"
;8��=Q}�^'$&�HV)���eF]d�>��������Zm�*��B��~��F�Y�9a{~��Z�������P y��8���(��MPg�D�NC>j�80�.�@cQ�^���'����4�Z,�
*�kѥ�օ���9>_�\������m*����j ��m�c��#Ǐ4w��?����N˴4q��o�\�E�Wll�jG?	7�w�"Y�w��Qَ�I�[�f\f�Ϟi�=��g�u㐈���{���f65�~�	;<�V���w��������d[&Z�ߐƔQU��4#�(-��C���4�$��j��B�Y�8���4�� s�����+o��~��W:?t�������i>�&�c�/����e?Wϴ��~=�ǝ��NbS�G����g,�~1�v���H�ڡ� �vMG`�[)����q�+��7�����Nk:��j0�5����e�G\��Z�h,ߒt��]�(F��"�y��q��V��L' �!��d�.�����3K��� 3� k�%ȣ����ꉛ<��Ȓ�⊝��>�IRO�r�<g#c�-?��P4���Y���M�9������]��l\�Ÿ,��V�x�zHL�E^�~+����B,b#䌃&�1��Y�b�E�w��y������rLxU�%k�O��*�뒄�'�MfJ��h��Or|����Y��m	^��Y����Lu8��)q3}\ߦ[V���Þ�<����a�W�5�f�sVZ�$��ݹ�CZ��w(���W1������x� ��7AT�rlT����0�q��D�P"|u�~
P�ʻ@�6�q��o��J�H��p���k�C�v���5 ���s⢤@��)\��u-���O��H�[��SϠ�Zr�!u���xH��AV	^G����!j�ԃ(!C��l����w���:��o�y s�u}���\Hһ� Qi����sѵ��y�3���)^�g�o�/�B��4�W]�����$@N[�DsW�"�
CZ��r� $)��L�<R܊���~fƴ��AK��������:��[�}��`~�4����/s��-�����40y���W������2|���Uꬌ�G�:H]$G9�Y	���W(6����59�������G����j r��a�9&�_��W�-p���-	 ���X��[����7�/QZ�����%}F�����UW���Ţ�@uڤ��v�I�^q����V-�Br����F^`l8?����(e^4��d꙼���[�h�ɡ\�����y��]"|W+����c]�8�O[J��K_�梿��߬�?�BS����mty�AR���!�d���p*���0��-I�o��uJ!�0g��n�?-
Oz 9V}zy�CD`'��ܹ�@D/�����&�u������Q�]
Z�8��#%���ܬC�VI
$n�`U�X6�M���Qx��R�ʗL�d�̻��+=�񰳤?5��K=%����IR�Q
� *W�U�>%Ѣ!��%w�)�-З2O����]00ϕ�����P8��F?�EDEX��\�>S�+���wq�^���{�pё���٠��'�S���IĞJ��ZȜ_ix������b`���Jv>:R����P�axUJ��Gc��H�4�hiE/W�������C�[�25=A9G�^BF��/~GC���c��l[����r�|`H|y�c��h���T�ʹK�:8cM�;���5)��q%�9���3b��y��y����O�2�<�6�������=�{i���f�Thm!�9ou#�Kv�E;XQ�K�aEw�nS�K��Bv7��[��6o��.{	]L���<�|Ѳ�[��)D����뷣�	��Mn���n%���*���~%gQ��},'rƶ4S.���Y�͞�[񳙗hHV+Dh�ЫΡ���x'��(��.�'��Or��a@�[�NRiI�aJ��tȂʓ����;A�<��^+�1��A�[� ���H��#D�|��%�/Cl���.�� 
�n�5���{+!�����&mA�~����
��M���a��A�o-<۹J-�
�YҖ�� ��zg%�TAp�����s'x�R<h�5l��N�3H�L���Td�R�4���˛�J��o���`��V�;E�;^�b�������ؑ���-�/"�ɱ<[��v����I�8� 1�[�&a���xS���M�ŉ��OG��TiE?!1���x���0���E�j���nR�RC35J��� �Ț�-d��;�>z���~S��c�}r�iu>a?����vo�&j��~��AÖ<W��s�_4�S��6�q���n�L��H�^V�jq�#?ycW���MƵ6T"�:,N<�^~]�e���z�J�����A[ ��لqozt�W{�_@\ ��i�^Юn��N���dwoA�����8K����&d5�Jz�oLk��F�HS�zr4����4�m��4)��Z�}r��'ѱ����_'T�^�YO�ep6��r��{��Q����|�H�NE�P��q,5]|�娂��I��8<��x�X��Q�%c=���� ���h�le=�n�S���iEp�y��p�?G�yZ���[63�vy��M;�`�z��V�d�S$Ym^�W�.����AZb�;�h�k��Ԡ��M��O���L�n	��#\ӭg�t��$�����97��Pxę"�o��v�+?� Ь*1���tYZ^���
�]�����;u�Ǯ��`aAЇ��kz��.�+2���ӄ��޻
�G�9͠��8���7��|�F���QO�0�t=��ס4��.���x����]W
�%1<��F���=��ϋ�y���5�7������+ZS=���h�X�F�<<�%��f���[w-������K�Q(���e�NK���h�u�O��G�Ztg�-R�,R�Ń���ɴ�ʜ��Jw���bsީ*цN0��/K�kN}�
��l>�Sgm�т.u�`��5�W�BM7���Փ�|n�,YZ�&��8:r�qpbIX��V��F���6��O�z;+}"��ž���	ͅ���LћV��@wu:�$�4���[��}�f�D�w��ꆖ���zF'v=7� ��e^��)A�uX�v]��Y9�ڼ�� -�t������sK竬m�aq5놪V� 6� �2b��RaI:��_o_�jW.��1�A���U�Q8�*�P��Gw���[�����w��<����)ƉWJ0k�ׯ���{IB�g� ��hgQDY�13�A����uʛ�X�e�O���W�����8�F��c(���h/g5��e����3e�H@�Tcҧ���ע�����`�JV"V��E���9���>X�Y�4S}�A�0�_h���1�)��t�[:�o�K�)�bp��&2�g|n\�VW��b���B'�KX[{�Y?t��`��zǵm���|<��Ӓ5�r/#��6Я�e�!xÕ���x�	cFef�?_�y�u��?��O�l�#�-e��� s�Џ�v��=ז�Q����T���]���H]�,�Ǯ~?���>d��
J��\�o~��hp'L
W�
��[ ��v�ť�"S��\ -�9��� �N�^ςRn��3Y��`�02�`ba���,�1��V�����к�7m%ɹ�Ի�w߱��xH�����S����"_!�)�z%�5�#���Y��l�=�3�nz�jL� D�}\X�ˌ{Y�D�+����h��8Fy��������'��լ�g4Xs�������c2�����b����z�V��@�T�?�LW�´���v/y<���G�y�=\����\�,VC���J*\���[r碫�O��"���^B��t��D"��9Ok���ɟ%V�{�*?|}�P��;���;v'���
��T��_p0GvI�z�8N]d4����뎶�J=��66j<���:.�]�]�5�8#F"M.>� *�,L�7�;FԸ��=�&$���&a�9:�;��h&��%]��B����$$����jv\��F�J'��"Ύ�����%��k�uo�)���c�g9��p׀�S�z8e�Q4l�z��>�|���pl���B�� g��i�K�Z�%�у���y�zj0����;��͇�F��u|� -�΢m�c�ݬc�Aү��5-!������Y��lӚ}��{�aE�BC��ۯ�`Z�g�ou�+�=g9v��<V�l�Eg\�ܟ������g�q��X%=P.���_����o�`�+��Ɩ�%�ሥ��F6������V[��l��nI.T��2R��U�^�eObZ���N�|�5��e���i�m��W�g�W0�*�¥x���֎o�����NY���ك/�`@>c�uc��-x|Z�F{TX��VeS�.p.���R��}0��H�L�	���n ǌ�x`�ap����%�=x]�ٕ L�x:}�+a��4m5ˢ�ÓV�=��P���
�bS�]
X�DnU�0���9�r�L����Fol<�d�[<J!��}�I��0�����g��i�{}����ϵ� �4s ��~#x�|B��v�}�����8��#�k��	�%�Fy�j�-R��T��&�KZ�t��0�����P"��kTi0ź�Ǉ8��R1�� @$�[�n8����_�C��A5g��9d�X�z�E�P�!!�{3&&p;G���.q��̑��,��q���r��R�8{b��!DȍH�i���n���#�D��L#������k)�ȵ�����#Yt�6߈�<tH4�K�ƥY��cv����vy27���\�B�&G�N$���i�/-���u��{��U�~]���U�YYl[�t��Z��|n��2u��n.�p=�6u�tR��b�ݐ��~9���B�XB���l˕
��c�4�8~;gT�S�ծ��V﷐����7�녵��F?�Bc�2=N�s��&kv6(�Nɴ���>q}����Jf�:~R�D��IX*�����/��j������f"�J8p2�\q�l��)��D��;HÌ��@��9�f�0�;`֨��o�ʁ�~"c]|��\[9��U�B��v�GǪw��?
���3�or�!L}��X"᷺�
��ȑ�ᑽ�x\��N.����fU�(;�u�M�5��ɱ"O� ��� �nHW�5d		�M�)ROC��H�k=�N]l� *���!�f�+��P>Z����RyGj۳ż��GL)'���=�{т?�ڜf�{霛y#۟�Ei�m�Y��-x���	��K���l���I;���F�;6�����������Sw[���E�X+��I_�{
״����e�:
_gAa�ʴ����^�ŅC
��;�7������� �?@�r!�]?}Ü���Z��{�sӖYJ$����R����l%���6�T�o��������#��n2���C��X�U���w�A�@�k`ےі�3�����8�:[�~��5#���j1�@�y2����f��<:���:!���K��=�L��t�$��_�;���S��\�w
��mh�h'���k@K�
y猲k{��-R�0�L#���
�RT��إ����Zx1���W���0�s��{��`h��G�V���� �����K#F����}�d"���Ƿ��+�#5�jp�FO��ij�D?#�I�TZjDmӏ雛љ7.OsR�2��36ZN;���������4|���Ѓ�T	e��`a�OX%�%{!��H���ݘ�VP 4�C4*b
pvv��!�6��HJ�k�ކ۷�a������.n��<�LMp b"���xI�4jn5|	g�)����W;û�� ��nf���Z�JZ=��� ��Ot��C	#�Y +� ˨:WA�\ �)1��ZЊL�;�[P��/"���,ū묽��Yo�F2�?��6���ـlސ��t��M�:�'���y�'Q����z�X�]׶���� ��*�����S�KN� 7�'u�{H�֪<��*sXf!mw�M��{�������[]o���ĩ�d�5o#�!��4W7,�s=~c����a��$�2[�]�~�Gn$Y�wi[o��T<�ʵ2'��h��ZW����\���.�XW��+RG�Sʾj��Y��'`����e
MS	���Q�'�i��S�Ê�X�L#�yg��(n,O�V��(X�X��F�M����JRd[�E�i�V�i<�>�8�Cz^g���ml��ث�jm�Omtp���
=�=��h��C�m�鐔�C?�]`�> $e� ��*��x��Ar�W�j*�."=�k��Gg�#U��
a��Rn������YH��M��2�m�|����E�Ғ�7�V�ңL�@�}���O� ��q+�ΣUݯ�L¦��{[�}��U�n���}�Z�s�l�t�x�yb"{.쬵�Sʋ�]��I���0
��#�����̡�q�<!F5��8����AH�֞�ۤ,ިiX��Qy�v�m6��̀:#�l��L����$��q�9��
�ء��EZQx�<c�L�g��=D����|�l�3�R��H&,�vP��U�#ױxU��݅�9�%� �f5P��p�B�\b�>�@�cɩ�X;<��w*b�����,��P�_�D�hU^4�I�y��F۱ǣ�='�%��Z�m��K������ÝЊ�C�ԟK�Y�<����艴 ��Ⱦs��D�W�d	�#����Ǿ
ܫ)Xs=�8����J��9*8��M�D��DB�*Q��f���?�˜A�eg~�4~�Rӯ� ��b��������]����o�g ���P����L�kX)�Bs��ҖM�@�o�=�h*�x��Bce�ύ�j�-ݿ���e��LU���ڢ;��������v@�cLܜ��v�S=�������f3����:m�{ߨ^ƣ�0\3�dZ��<\t�v���p/�"��P&ɘHH�s$Ij��5��9Ue(C��kM ��paVA�g�)�����w�و�+R>Mfl���NHO����v	I�n�J���+z9������~�����3�%��,�O֚��ñ���g��L�>��]5;�`җoJ����h��ҩ�Vk��D�L�P7�{ϋ�i�n���t�P��ί��?�+�������h߳'G�V)}���?���'-JW���yDR�7�ɦU��˰dbd�����#�8?�-�}.3�y3�m��d�s!�~�6!�{ϼ<*���H�r폆{���P�~��3����"����H��yՎ=}Լ� O���YB�����ϸ�&�g�(\�����6?O&�apMM�*|�1_.>(h4~��0@2r��l��h� ���ǹ��^M��`�a�ڜUv����{]H��(ה"�:w̲b��~�уmD��&�]�/���_�c��{?����:p�嫻`��~�t��SCv�"Ay��n�CA�q	c��K�ʍ�w�������B-�sI�qij��!�AZY��ݼj��܍<���XL�}4�i��G�\�F*ٚ�r��)�Еv�HW��t�(Yiw7�]����V�l^ʼ�kh����sN.
��d�u;��:����a�_M��mH���w��I)�����Yx�#��!��x!��������Oc֣{���E<��F/��^f��т��nU<iKyZF�w,�.ey_D��<�<u�0��o���b���s��Q�;���j^D�v��/�78)`�� ��h�ŏ�܍5��}4mq�TFg����1lfI52��]���J<�]O�h�X�B=�5ʪEx���<c��Y��;�6O&<����-��d��P���[c��:Yͽ�b$�z ��'�&��z�
q�����֭/	�78x�p��5*H8;4yX!���H�|X�}�cg��&g=
T7�1;�)>ݰT�\�I1��hZ Hh:ހ��a�m�l�8K#�p�x��:���C�Uy�J�� ��`���O�ΣfF�E7��NᛦW�
�~v7Q��G�LM��B��}{���U���2z�u� ?`��Og���gp��M��ώ��Eg*u0����a��(���\�u�	���	x#v�;g.:&�����a�03"���BX�����S$�F��k������-�cF�N�C��5Doy=?}������RRi��Y�Z�u� 	B��� םa@�Ml�n�LxJ�1m9�^TQp<ޢ+��jcm���`1A=��?�y�VQ��|�3��|^`��}�Td���:]&0���W�
�h C��ib�9F��X�7�¿�_(�F�=۰�[R��L;�ڼ�nC�wo�#��#��ݴ6��f���QN��M��zr��V�:��)��!�ÍD-������$�6�/�$�K<�l���:��[,���nz�~��i��Er�R�b�z��I�sFٮ�54��2���8�#�[��K	��M��%��=�b|�z�-�J�1Q��F��=U[v�8��9�zY�����t��V`/�^�W��7��ӏ&����k7i��>�T�?�I3k�^�p*���+(�$=g��9Y���c=��~�[z�U��x�d�I2��B�~��y��匓M�GFA`d.��t��:�
�s��k���v��gA�Iw��M����z��w�ܴ������'>W���5�kA�NĲ�{؈�v��c����]Gm�BE���.	�B��,Q}��ܽT>*r�BǨ!��7��u��{���'s�A<Gn�״�R��D���_L�G��y�;	eD��)��uB+1
����CcR����O�PK�7L�k��Db��� ���  H �	��ms�i+B�Sܺ�G4�Z��^Kh��D{����G�Ʋ�ݙ�ŭ3:���Y�'��Ì�`zA �>rsR,�[��������U�C�͡��i���M⟓�Ք4��X�f┻��?l�R`4�C�l12��"4�g�� �H�Yz|��k��zۮV���U�B�/�-��jPa�Ң��:�4�@��?�3C1�}�ԛlnT�L���$�|�c�ѱ��Ħ��(��
ۭVa�ed>K�O�}|���]N.n�π���^�u��m'_�@æv$�~6K�W�|؄�k���=zm�0��e�5�I)z��>]�B<u�5>g%��k.O׫��<��h\�Vn[$�\��ӣ3zO��O9�\H^n<0�����
Z�	Z�d�����o��-�py���7'q����'�O$K�RS�對�Z�0zP����Ąx͗�����5v����t���f}9F��p�t�
�)d�s���t��tqW:�g��pl����B����e|LMH��N9�1���Xd�B�l���x�Y��1G\�� �꿚��R��&���G\~}���P�\�3�@%���l�����p0�t���hZǗ�����G8b��C<�0>0�'�k��Y��'�CU�Qa��O>��|����o���M=l:^���g|M�!*��6�9��OI�%������
�?cqȐ(������o���d]o<�h��V���6=�X�1�>6^��&�{������i�*	��T�`]������������}̞���eR-�@�Y&C�{v�+�_�\#��P�Xji��m��W�V+s�6r^sW.:�kN�<��z6h�o��D�}�X�W�,�ƥfz�]�;�t)��rI�!��DI�}y�m���H(�W�{85���M�kw����=[�������w�t�dI�517��*T�!��&E��O
�Oi�d�d��������D1_ƙ���w�~"�@�y<_�w�	lw��C�yko��ޑ����o3��>��G�G=�Q�q������i�V-|�Y��Y�(ՠ�QE�8�L��f��j��zy�5������'|�)����Mv�~�C�x˒#6Z���A(�ۿ���nYs:Ʒ?�<��=�������?�::�@��Q����D�r(ֆ3b	�H�m����-i��yտ��z��ҳ�[C�f˚�3h�I� ���)��@b\P�1&�$�V��{�v���S��g/·���'��@�C/����������n&�Z�Ów.=��>g��@�R��E]��n�(#N�=' �𦇪-�3�U���ߗ��E��@w|���2���y
��|�qwF�hݨN�����OR۹L��o?J3�h���r����}�j�z��QW�}bF20������/��jI}m;�s ���z��8�����񷕞r�|�#3�0�X���@A��`I�kQL�-�����q��FPqZ~"JUGm��R���x��G��������T�=U��o�E�~�]{%�c0�C2K�7�C��=���;r����[��p��_Р�F�ƒ�o���6�-�N߼������N	�%����5���bBˤ-��.�m��_�RM��1����r[ۆ-���RJ�U�*f;�_,��7ͼr��� �i�nON��t;�Ϙ��f+��3���|�_�2����D��D��
K�� Ōg�Mѩ/�ZOs��|+����cy[H��|�����'+g�:{��!�{���w��̧�O�ZV�8%o�q�B8� �D?����l�(�K"œ���(d� �s��4zT��v�b��CPm��9.�:��ox0��u�F�+��/��׺�<�e��g�'��7�OE�	�u�>�.��\Ԝ�<[�c�ƺ�P���0N����7�2�e6{�m�����@�� ���2��t�+�\S6���E�����g�C�9�\���!ӭ��.R�Q�Ё�{�\��C���$��y��b$���>�y
C% �̩��8�g/{��+޽��m�a¯j��{�O����2D�21�p��|R�j�C������V�\
�ot�98��e �]�puC��#s�`���
*�l����r>D��͆ �f��P�\��&�k��&��]zb(�wzXp����Aْ�,���$#�*Z��B����7]t�Ǹj>Z��[�sJa���-��9Gp���uWC9�+��R¯^
5NJ@��7o�A	�n`�e����֣y�N�<��=�����菓�8#GB;��]k��G��̟�9���87R����'��Cn�����Yʀ@�X~.b����q_�}Jk���QKs!gG���2�b���D�����	���.�h�xo��s���]�u�@k�h��t�B��ѩP���WX;Q��Ȓ)I���9#yɴ�mka�us�d�ϧ���`�2-�K�'��N����T<ש����H��M�:�?&�z��|��ם�4�S��d~���d��L�I�]���V�U�9?�Cuk�Qk���b�c�%��o6W�J�o�3yC�^��Wn��^�̘�Cfq����5�}&ts�S�}��Q��9~�|��Єt�@G�ĥ��5O���,~	CUs1[9�������C�/��?���GݍV�������GK*`5]�#=_˺M���kY�\����tN���	�m
�\�x,V(����~�}#j�t�q�@C[nM"NoG���֔&q(�q�ܹ
����"�_����۸%��wfvT�[���űl�/.>���Y �u�m�����뇃�G���p7�Oe����AG�z�w�s�j�w�5?�y:� �;E]���Q����S������E�W������}]#G�ͦc%���rw�h�����a�3�S��E�[,%mݟ��,|�fE�k�h	۵;	�z���S/�W���1���s���Q)�|,5y� �E������я<[j�p˯��oOܶ���q���EDAX7N�ن�]�tuR�qi%\R8�np{W�b�Z�"�oYA�D��,J���+��;�)�F>+�&��_��s�H�w��.�N�A�}��mF���������[�UX��D���w\g�q����L���ܜ���d␳�Z��Ā	c�qϟ���o�U}������x9w���dl�h�U��z096����/+b��������4�~�)�T9:�eOSe�Pz��v:��m*@`�����(���� /*�7�I�[)��D��C"��l���j�^�����S뭐V��3���<X�xO�I�I ���k�E�֡S{���6��;�*8�?PG�>>-°��1O8�s�Ō�lG�w�XJ�.���$�I����m`US�E��M��i�@u�o]j̰>-�'����&mMu�?�VF*�գ���黺�o�s��Z����,G��2k��B�t�t����V���؝:y;���:�nd��P	%��Q������V��~;&� ���FI�����!�` �Be�[Ԕ�h�U��q��6PeF��!L���A��S7gf�H��x���?�j܈���]����_�/#wWz�t=�5]82��>n��?���L7L�ֱT�(O�]1�
/�ᦳ	��x��Y�!yV�Y/
p1�[fs����>}���s\���g���	���p/�_���*��F�AI��D��d5DְJR����:�8�Mw���/����*���e8��4��]:�1T�(�ʿ ��1�Qȡgp+F[�"��,��b� �+(�8����#ݶ�_-�e�'�j��qRE2|k��?��F���<*�j�M7�+�����z/�����NO=
1�?Y��qf�H�2��i�lRca?')�t76�\�ls���Oυ��Ѯ��4���͏)T�..z�H����W��".k����|�RSdr+ǘ���sQ�$G�B}Xtr8[#+���!Q1վc�bbk��ʫ���ӅsNg��������.�2���w�*�K�(�*�W���_��d�RF��by̵S���VX�Ge~�<|�]�xe��E2�C{�'s2�#��@���S���ja���ԑÉ��J;�?���w��g'χ�Y�ֲ���g�c�f�0Q�3�������E�V���
,q	�% ��H\;MK�:����N�|�n��D۱��;̡A[\pbU��c�]	��z����R���ޓײ�"&��K�=��g���I�4.F���$D'�</m8�k�t�i��9?��p���P6��6���%����D���f����z��֌�Q��]"Έ�ݵ/���&[���ߚF�nG5���sd�ь��z`���՜0m�E�֍?ht(Tj|�b�6�d�y������2���G݊����d��L2���?1:�#�S�k�df��m2ۛ,�#C��>�f���[i�fO�m���@�>����>���B�{�b����U}߅�E>@[.�B�Ib3��:q��'��a�fb~xjV�Z��\�T<�ΐ��a��Zl?�2O�����'�-��r��{2���>T��>|�?�¹�q6}���|. Q��P.Hn&��!�輵��f/ަ&�2P�����k��ri�ގW�D���0s+sbSr�ϔLG�O�J�8A�Q2K ~gɡr�Vۼ�	��t)�����A�j$~��#w E���{�aX;�QZ�Aڀj"��?I����Q
�Ԍ�^�hi�;��Q?M���ͪ�^iڎ�6꾝�ѤΪ4r���ic�HY�:����������x&��\�ˠ��{��z.'d��묛�f��lZ6rQ���^:�(0�O�H�	Ӻ񷽦A�$�Ug�	���KWm��`vx���z�	7x�N�}besƘ���:��M�2T�0����k�7SB���e��]$�ƶG�Ƞ2M�dR7p۟�	�G�u|TK��e�ں]�L�2�
HNSp�ۈ���+���]�U���4�tm\�DO�E�;{��@3�B<��U[7�G١�E��nTj�Tk:[g�v0Q10�jO��t΁ɼ�V82�V��O�9rk��5/PN�6�/y�N�'�*1՚�������r��Q��ɡ��e���|�֫`y���uʵ�@�T,���<�@Nt�9,��K�"{1Lrhv����h6K�.�0�Mrdq�)�p$�M2G���f�>e�Rk��/D6���Mʱ�ǟ��:�%���B���I�4�)��gQ�Ć�B'���ozKН?
P�(�_�6��Sg�L�g)=�e<�����9u�ΰSK������<������v�z2N��"�>�~���`+��5�7�ă��">J��a�#KȈ�SN�`�����1G�8���"�ƫ�Ġ�x��J���ѷ���D:�K�n7��T?먛͏r9_���b w�w5��Y��Z	�*�/�=�7._�F}��Q��]#��@��+B�d���T�������Q(�oC������K�/�柕n��Ҟ�׹����r�eS�?E�{��VH�JY�>�k��O��#��O!�ՙ�Q'���W�������tc	-�� }nz�2�9Z�����Y�Q�k��\��A���c�n8֡*������ק\��mv�r����R�X����y�_۶��Xt3��e�5i��>[B�8g���=��$���:&�s�y������>Rf�q>n׺���v4鹜�qry�=?w��n3����C���_A��?���? Q�ɪ�6a�;��j`�Ϲ���i���~3m�wb %��:�L�L���
�}��A��1�����K�C`9�O��o�@7�����=
o7��a� _P)��\���r xܿ Q"�$��>n��Sm�I��U_rf�8���{^�IJ�G繜��9�C�t-�$҅��b����W��A)5����(�!Q��?T�2��^<���#�D���=Sʻ9��m
U������K��f�S�dO̎^x>bKA&��X��O��b��`D�@G�M����{�FɌ�L? ���7,�a��6Cg�A���(Ec֍w',k�՟�,;��Wl����[tW+ �O���3љ�w���U��F���)]�]�8<��&��/���@e7�I�����Z�Zk{��v6�E���q��|�h�h����ģ��U2 �MI�:XE'�+����_�)
��aASi1�;�K+K�sy��g0�L��6ѫ�����3;h,�j>��D��<E�{�UD����q�4&�� ��l�}<���#�&q/��>ř���P
�ܩ�'Ğ�I�+6@�W[b|�FR������Z�>h��q�g�񼯇�ߝ�����b��Ɯ�^uݔ�/����g�Yb�%E^���:�R�-J��
X���Rn}��`���oC��9��ʧlE���d��K�O}��6Q�r\�9�7�+��P��포�B�ܯ���N�X��	����l�G���P(����l�J�����!�l9���H���*�\>{k�q��H��}AK��"��r+��?�Ky1������W���+XAbDc�f�#���/��J�[�bu��y�G1i�J)���
�yε7�wВL��2�����֤H���Z\Pbm�ë��-�5n��+��U)��-��6'�㐸T�Z�M�]Ƙ�_+��n|�a_��V%���6W�x!�n�*B��J��g,l��Ѡ)�k}�wCM�Cdq���Й�1�w�\|���$E��џ>9��/:8r#7P�ę�{v��f+'.���1H<��'���2g#֖�R���.��J�M�yf��>�DaASN�k�`80����L4����c���b��R�(-o�p_� ~ۙ�hL�+�g��S`������E߾�c���Im�vL(�`��{���81�N4��0"�lJp]�.!���l[��T:mE��M0`�5�\�&��mY�f��������ʡ�7�L�ۣH�:9#6��?�X"p����r������DG�cR��Vdis$��]�&*B��N�ɨ����h��K��ą�i��K��ˏ�5K��!d�e��;���=�p	Y׬UZ:�����Z �Ҧx�ꭅ8c��:#V� ��eA�y����W�k��A�;���F��'@ܦW�Jؗ�u��O&B�:��t00R?KA��6�j������!x�u���d�	�Έ�%c��d���Ʉa�~�4gjB>$J^+�x�'?H����%�C��A�ߕ��Lx���W=�_Ģ������!��\�G)"���s�T�s�����2,���PH�5$��)��4e�?����R�.W�q�j૗�~�]q�?�;B�|_��῜�}h���R�3b�̺A�|�e�+�4@�Z-��bD]b�I�������p��E�a�%�v���QM_�@�]�7���1�B����QN/�����D�.EZ��X�X^�!8\,x���|��S�<� h�G��Y+j�����|��������3�� �
�Ɗco�(f�����`K������"����l�M	�2���)��'�=�&��Jԓ#bC^*&oO �>�W��X��\��U�k?��Ά��Lř�������K]&�9R-С�&!��_���	��#�L��s��b�����lCM���%��Fd%�v,���nT+*��4{	���W#N0�>�'ę�PQzK��|gTS�ҿ�r<�*�(��4!��t� ]��@h���j����J(J=�H�R��{'t�#�����?�k�_�e��v���<�L��<��|M֡�XV�����<A��6��|�D�U���i��iH��[����-�3H����ne\��/E\�e$����?��_��}|U��v6l�VH`�5�ז1�Ӧ�ݒ�j��6�QB|�� � L.�,S#��Q�v`w!�ZI��5��U4=�&���c��J�~$k���Ti���@K���~��O�{e��sR�-��(���-�$Gzk������^�iO�;�)��DR\i]��`f���,EB��'��g�=�Uh�����V��SQ9����y�X��@,�iD: �$p�����*0E�����j�(��h0oq�2Ъ�9�����qcrw6��9�L7�&�9\���]�������(# 侽Z׫FI��9�����7?�z֏fx�֝ �0��y �����)v-np�?�yGJ�i̒�=���`���!1a7X�F�í��*���>v�'$Bs�� �����$F���-/z�THl+���ϭ�T�N�@��&�\b�-����_6G�D���=>���)�5u�_9�#>d���0A���(�/�^���j���y[�%pH��y�Y�GR� B�{�,?V��3�C��X׼�P�r c�q8ޝ������(kJ����i��VHI������hw�9�Mb�>��l�jN�Cg[�`���$��\�J�3[����D)�!�ͳ��u�����fq���1+q����8�EN$>��<�ڞ� �u��{L�_=�-G��G�F�J��iih ��7��w�
ĥ��6K���~��Y-���ě�3,1|�w��$��*qI��;�&[��j(��H�y�9S$i�S��� w7P�Ա2��&'�����}�ei�q���w�W��{Vlڃ��Hb�z��]<r�D��H����; z]�����v�>L�%:f�6�`�kޕd=1l3U�����F���9P��Ʌ��(>G�ˉ�_��+6�"*�d.S�{Z�c?��_!�,x�绶��=�hH�bJ�I��/b�����5brʯ_��R�_AN*��Ai9ֹ���x���V�ON�;������~
��l�_��=�{�׊�J/c̸�[���Q�@Y���v�(m�ܴ�RI&<|3u�2�;c?Ѝ�Ş<��~>lU����Á٣"^�Ie�9�
lC������P�#L���*�s���O�^�-}�D��H�D��S�fyhM��v#�͙��e[���h6�j�N@(�e?�?���3�;���wF1�40_\sV�joe���׉ ���}��9�{���Y�~��I^�2���/��|+�����j����ҙ��w^�1ryO���b�]Ӵb~{�|�yƺ��&�l͹����.�q����6�`<�A,����B7�$�4�1DV�H�S[�)��(}M����f_.sq���Щ�K�6���;*�]ju�'�������0&ѓ6�g��?��ҵ֍I��k���b���j��9H�0��?�}*
#�Easn&��E�'k�m��vJ�/��yu���R-L|��%JK��h�'�3L�j��:����'�P�ӧ)�p��i��ީ�%o}2�t�|>e���:h�8u�e�O��בݩ�W%~��_ݵ}gl�9�@���,V�wVP�ӌ��B���Qߟ�sA�	�3V
�}T؋L�}��H���V�5g��5i��Իb��\D�<!�ǌ�.����Q��n�k�>�_>�u+ɢ���&z�����׾4�Go�p�S��+`��j{v�FoEx�
J���a���1��ԊL���!hk���m��޼���g�e��Q����齻���%d��^�	zb��fb���_�G�s>p
�$����ck��ɬm��ú
WV��
�&G��"2O�T1~JOfW5M��ΊSc*@O��7����bؓl�12<Ŏ�0����!O%|�Q3���7ν]N~�4r�CԄ
�(���<�
��!ZI�7����E�s
�Д�ɮ/�5Cc����<DAN�:��U$���B^��	�����9ܚ�����[�1!]�A5˝�-�Ԫ���!���<)�j��2�K9�q][��ػ�+�K>s��ïK�C!G��.��db�@��#+A<֨�[������s8l�,7|��p�͛�:���񮢼��Rc;�Q g-VO���	g��ᚾl@�ȎSg�N���qP����`�-�U2(��Bxn���^�ZB���w=�I�t����8(��F�Galu�Y��\�҅ ��bP�E.��3���?.[Ⱦ��h�n��E(��6�{�U3��V���:F���U���L^���;�����>"�xD$�݈�Z�gD����n�l�p[:J����у�^���*E徕�//:s�;HK��&���ļ���yy������y�m�/��Χ�PC[Wb�猯u������H�#�g�T�y�E�Y�ce��<>W��:��5�Y�қ�"_	�����g����n����8�n�nK󕼛��*x��Ss۝ �~n!Bz�מ�6��-f[����[^�s�� eM��MǼ:��r=��@��F��s�~���j2廬�M�7��E�|&x]]'V^�����`v�>�B���I���V)�����2���I6f�l4=g��7*4a�� �>*~⺼�H�pIM6�-iFm3�����]0[��).pA�u_GAAM��P&©�T||�kH-4=�:NE��8�H
296����Z=~����^7-��u�~>����m�ys[�� ��|2���E��+O��kq㥵����b�N�V_�&�˷�r�˴S֬��ļ��ng�����WE=�\�rݼ���6�ƻX���=�|��#���K�Yd~S���{[fl��AȤi��;4��� ���Ҋ�.����Y��-�f!�e�z��������Dw��+�V�6!�>�|��xW�ڞ���B�aޜ�a=&fEҾ%�w��H�N\�
q)�s83��U���<ٵz&���:�*&C� ��I��T���wW��t8"$DY69|+M��w�辯���?7q���cZB� �ķ���F	���᧪������x�EQ]ѓMz��U)爛t�B�6N?A�ֽL�`C���w�_-��EP�3E��N�]M�H�q"D����HI{��3w�@m���jF�$�6�ZJ �B�yx��-�Vi]�O�<S�~�k��]�.�I�+���e�_v�����z��f�Q&��{(뉡p�+�s�X�����H��B����j�"5��|Zk��$�=����+=��?`4l�k��"����=3Qx4�ܘ;��Fn&]f�V���Q/D��z~գl�S]ct��ڠ~:�h�s�l�ב�Mzѵ��W<HSUiW���.��aH��O&�0U߸qRk�SM&�i-�yxńY6��˜O�5!�Y���<�(����E-��=�~��ˡ�j��a�5�����ƩU ����U�:C}vaf�Z����U�e����(�TWTjm�*���"
j]kڐ#B�Ć�V3k�^��U��wbv[�R���UҦ���b^!܄�xL)7=��<Q`!��9�9���g���&��ز���u����(l~�I��Oj:�*q�-C�x��[����d�ƅ/o�sh�
��m�C��^*���yB�b�ʑ��ؼ�`��B�\���?*��8�o�:�vU���gy�)����x"ڋ!Mc$���.��V����<�v2�mF	p�9�'�f����э,�vj
W�����5�6*�����ٻ^D�ϢۣD���&S�Pz�)vz�dy==�����2�a�5����M�:�������p���Xt6N�3G�0������c�>!�UI)z�X�~��YNs!���86�]����$UtK��3���*������6�\���+`�xU3�UQ��#=->FnU͒i�I��z�c&�҂�i=	�[�����i�ڿO�f]Ii=K1�[�D�A2b���S�]���"��
f��a�����Fs&��E�9�/�!��]&�����d�J�=����V�����>G������r1P�E�x�A��za�����(f���0*�F0^��c������l�sE�Rm�������Z�ΈL� 0�e���!�*�>�&�N�BG3#߉:���F�4�ÖP>a;�L~iɔ��u�lhk�UtWN]jdcFsT�̚e��`٧
�i��}�Hk'�'�v�)�0o��=���ꅽ� �; �5��9A%�-�3��C��!��OMY���)��՘�oÄ'M1d���j�>0�vǡ�FV����'JJ�7^�d�K��Y��Ĳ�d~Ď���t��w)����e{�l�=���w��,D�N]��V�A����Co&~2�����d�%��r%]�9�_A��RZd�yv�L�w�|Z�?��u��f�BP"(�Tm�6yS�s�,�t�!f�� �^���e.�5�ɰ�/B6MW�>#N�ڟϷ�Q��+�MNoǐ�<�p���;w)9�T��%�y�%�w�`j8c����Y�SȔI;�ku���ܪdh��'!�l�L{���F�:�<������4\��v��E,�;�݅�Cx�./�)��.�����iu�����i-6��j_�;n��g��_>re�oJX�K�27Z=�u����7m��ڊrǂ2[��:�p����id���@�D.)���o0��ZX��q� l�bTJxs5�FN�1D~;ʜ`��j_'!n��y����XH����2��qO�к;VD9��]{zr��z����T�:9����t��M�a�:����r&�I&����Q�����up�r�o̠;�x�茪r͢}���3t& �縶��Eܕ .RW�\j7#no�\a��v��E�v�yr,�˒.8��*_?ɬ��厏zsಭE�؛�ͳ���<\D�f"�<$~z��N���y��_��Ȅ��/'�
�X�ŝ��G���Ε�B7zu�����q���� ���AG=��`ŪƟN���Z}з&b�ѕ���[ZY�4� �i��Ui7��b��SB����\���O7��6�%JZܲ`�������ycD^X�90퓺%��3��@u{=4��*#3mְ>����Gh����)�Kq�f���ex��k@��r�5�2�~���"�eI���L�E	d�|#E�vee��&�����:aj�s��[q[����S^U���B�bEN�V4�v�a��\T]�3�L�߈/�jh4�H�Zv`�X�G����2�q�-��b���<����c�l��:.���L�h��N���K�x�!��2-�:P�)�$r�ʺ�)*q	�mu��XM@n0�2M��ݍK�)�\���f��y��{uP)�� +�{�d(�q�n�Y�BT�c�.�	��2<���lz�-P�}�Y�
,�P�p�j��q����	BH;�P�N_o+w��2��(�0`�d'�9�**���f�9�U�I0���@N9r��
�������7�l!6aT�9����Bp�ԟ�
@q�|�i�L�OL1Z����H��ۢ�r��3{���]��ʖƬ#��g&�DA�V+�"��{��1�	o�(_����T7����(��#���L�c����Π�O����:��hs�\+�jZS���u�����?9d/F��<�j��h���D��U�_kDܪ�v���L(E�o���5���֐�<����\�0��k_�ݔ~�o�df��|c*��&Ҵ/�t��'����+��9��:�'�eEy���.`���x;�F���0N�wI���1RW�c�W4,����	R����kgZ����D*ՙ��fɻ��c��GX:�^�͹���}BT:v���@Q��Z	��gdϣ�q�[�2����\��+�}���W�~�<j�*��N�$�@ԑo'y�!X�l�m��Ê�q�@2�5�"�����+\�E�9"�� _�#y�N�F&C��Gt}orѰ���D-�r���l��-���<����'=�P�eq���>�K\���(�S|A�7D����"$5h\�h�z>�N��?��S���ʂ��������^�$,K�Nȹ <��/Y�<˥�4r_tg��(&���I�0qd���"���i�
��g�{"�b�o���C.޷�~d��$��3����}`MG{ &�E�25����Ĉԭ��M l�����	Z�g��.ўrd�r�Ϩ�Ѻ�gg�ý#-�M����w<:�}��Q-�b\?���w�K���d��m�R��YJk(��e6��k����KxH܎^8{���3�[�i8��%×Ff꙲T"��x޺f��M���3@���$�����0h2]�G��+�#���a�v���I��Yқ���D�q��!S}'{x�ی��th�-*�ś�w����g��@�y��V��BL�e����.B ����V��"x��˜��] �+*'�a��M���*�����#���s�c�A���Ğ�~u���Y�ۼ�1��"��Q�ǂ*0�`�H6��%� ��𲎔�N�����?��ap���)��P�}��	����|-u�� ue�%��I1=j:8�~v���[�~d�T�*槣�c�EPO���X�L�n$�*4Z��o쳎o?
Q�T��|HA���ˍ�oϥ~�g�;��2q/�������\�_Ey�������P8�s�bɻ�ĝ�)�0&B(�E�z�ü+��-/?"#�E���[5a��%�}ZZ+ e"Doq�g���'Rm�U��*�����U�Gb$X	� �>�͔S;Y�`$��U祿��r <A�r2��u������#��̇9��W{���"�K`.Xfa[�U'ٜ��R��bh<��{���
R���*�* �L?>]��L:�Oy���Ot�^►1��b&(��*=G�6����2^~��s�VM������K�1�X�����|��0X��9�Ogz��@!ޜ�0IJ������M���u�}['h��ow&�_�hO�)��F�_�d��
r|k���O8ߪ����CF[�E�	�J���!��ʕ��Ǝ�/ɽ�������ukך�i���b,� ղ�pkB����?���x�tu�DЭW�PH��1'������S�R�$xxU(O|W�Ş��Db#i�����<���^,���Bo�"���HuA�2���#�i��F-YC�!���K}�.+A��P&¦�����)!'�ȡ>s�'9��ݥ�jNsO��QcC��5�eI�pO�◱�6���Q���`��	�rLaM���m�Ԁ��%��lw��Z��c)ϕ���y
L��h.7yz��Q*ɍ��S��Q��l�}�XIe��Y���ɩM ��i�e%�4�y�_���	r��LE��E��!j0���ɲ��)��S������`׆�Ǳ2ޥ������d�,��[��.�窘�J��7�߽���N#eRǢ��ɳ�8��>���	z�q0@}����j]��l�t>�)!_(VX	ݺv��V�4E[�N������3 �������$_�.��"j�����Jd6^��&�~�I���I8�H@$GT�&�bˆ�Id̲(6]����3m�[�,(,I4a������DT�k�?�\J���=��(�K%�:Y�H3�u2r}��h�׼
Q��u��m� �82"����%��L���%M�����Ċ8T��Ha}���[U�dX�>.�6+��'��tN�ʖO�ٰ�4��ƹ�NJsEa��/��~&��W�������L���zD�!�-i��1?�c7o�aR���:�SGg���pY��C+߰N��4���m����CZ'��N�I܏�_��4�i�C�"�a��Ä�$��Оqn���Yg�m��Z�̺�����'�{�V�+��f���{.M�7ʷ�G���135}^+��B�z��o��ڠ�Bo2g{�>jwb$��Q'�̐��p �7j��PX���[p��r�Aw�5e��M��W'���������b�1�n)^[F7��x ��:�����/iڰ������k�o����A-�\��Ǳ��؋�;�ͷ�pK��z/{wk�N!���V��Ҹ��u)i�x!m�������A_�F!s����?�?���_����G�/9S���ҭ'���8�������N���H1���?\��7�s?�$��_a�}T�����\b�l�255��7f��
`y^�N~��g#�m��r��|�;]mdĠ��myy�����NNN+�!��1��k+�h�����Pt��eT5���P�/���b���/��?�1m���������_�/���b���/���O���˿p��RCE[9�����PK   �e�X�/ w� /   images/b50388db-476c-4829-8b73-5cdf8357e0ac.png�y<�����]j+E
�.D$IY��P*B[�P�B��2�n���`�E��)�2e�,d2���yf��3ػ��s������������������^���s\RV��3��f۹�rj}&ì�y���tk��'���.o��7�o�:�e��p�������eu���v�v��v��6F</t����𺕑���IE��ه9'w�}�X��U�K���a�{��ʇ�B�8l~�`��8l-T�~��g.^}o��ņ����v�#5/\^�힜õ�l0o����B٘{�C3M�Q�ܓl5a��]����NѺ�f=��ec��ݨؽ�w6iN��W��q�����k������S�Ǡ(���ťKGvɧ�p+�+�0�����$���K`�"�#;540����	���L�L�>����$��P夒R��A���LWԔ��c+����L|�:60JZݎ������F��dj	�M�uWUU�xG�_���O��q�Qk�xKh����+>��o���&��!Y-^G�r�Y.ܛ ����t���Ա�,fxM���X�����E�v2n)?�����%M����]t�����Ӯi��}Lֹ�?�U�����8R�<(J�/a%��c���5eC������1�L���YB�0���O3>1�1ӧ���Ԕʼ��q}����CR�[�~��3z�_
_I؏�ܔ�"t2M�2Mp0Y��M�i��1YG	V��D��� ^���r�`���l�#ǫJ5,�Ϻk�l�Q�87.& �X��T�٣#�׋P�s�?�On�#�g�o�fE~ɼ��ȕ���(_��Gbn�S���)0�#�|���"��Qs��JL�W�*|ôjբM]Ej&"�Oz�@�����/�>]�=nO�"�8�Qb�u!�:�		������:��%�^C�	J�9��¼tO/8ZDm|4�`Q+:藞�����M�Ko-�2�����Xɍ�<�8ˁ�2m�!�c�.VVZ7��|Qz�=�Ȱ�^ ����䉧j���ev2ɰ1�و�3���䏡]NҐ�/b����	�9�����}0�3�!��Y�l~���\`�3�[K�I�T�!b�z��bfI�$7InWnn�LMU���{��9��G�Mp�k�#Q�+��vw\/����ݫ��(gKW�%���$�Q����3�^�(��a#����_x�U�/�-�>t�$�|'��vЀ%#�j,��5~�v�>��B��3Ž'mn4LNN�-dp�bm�
�Gt��
ŴT<�+=�&=�.���=.o�>���KPܫy�HiD�U~�*Lw;��e�`$�dYGb��u�&����ssVun0������Z���#4�#���L8�v�b#]k4f��&l�RO�o�fc�	�Lׂ]����
��DB/9Q�<w9�Iߋ�OX퐪�p�RA�̡I�7#�.B�}Oj��	5����}_�6�s���ˀ�	��H�C�eHZ/�i-Qwwg���)�a����>���S��s=���(؎,�I��q]�&Ԙ ׃ܯ����	���R;s�m2����V/�\�I嫜�R��<B����(T�R�H����w�Er��Ǐ�ISSsރ0��cpl����H�aaa�ei�X�;���ny��32jA2�'یB	�ܮ���#��wѓ�q~b*%) 6qu��Ȝ�����ZRZ�M�(��!�-d�
��7�Yyzݼ	�;�^׬X��+����N�\��	@gɄyV�T<�U�B����+��	��f4��Q�e~b ��H #"܇���3���'c��/�� ��Z��C��M+�v<�����҈	�ڵ��zl45��@�Q��aK�b?����J�����q-��F��}�ȵ�.��G�T�0��A�I�2v��^<Q��~�ToB�?a�6Cm��4�ε4g�~�7�3&�
�n&��Lǒ�i����g<WU���TJ�QFBfOW�v���s��?��a�FM�HoBdH/g$�z��� 8�DFҮ����ޡ�N�;Kn�K#��F����sc).ge�i"��p�ӓLL�SYg�:�.;,a�_�r``@8 �<}B���������S^��>W-^NN.��@ h'�j2S�3�����Jz�in�WǫDk�u��V�$Cr<�Eed����Ż@�-s�ª5ut|<<<��^�5�9:%Exqq��ڵ}�GTA���Ғ������-ۋ��D$%��g]�I0Z8�CEϚ3m�<�t[��M�&�%��pn^�����˗/{'*E��8�F�CCCof�gMqsG����]2oy�_AQ���Y������\�ˌ#E2�� �9G^4]� Z�������D;��e]���C�*T��xY'�&���Xơ�=��	���-��c-�<o�[w ��ٻo��Ԁ������C�x����c�2��!�ϤSK��66��W�[���W��L�;��pc-LX��v�[�$�Jb�Y���(5YΓ�� �kx#
Y˾���'ʂ��H�MF�I��@M�ԞX�H�'�*��ߟ��H���Η�Q:v�u9Ynݶm@Y��gA��j˰�^˳�$mznK^-�P[,��UMo��+�/�������hGy���U&^։���������+k�����3'=^��|�Ux�������zYio�O�5�*-.�˝����-�=��ڨ2Ⱦ{��Z�qt���h�%�5}��F^�N�`�UO�]O��
C&��9FR!D�/`����y,���Y������s���.��\Y��6C�{��VǺ�h�R�`�[!Q?�跷�͛7ӗ�:sb�u�O��=��̟�?M�vh:���:�/���`�w�u-��.��N��B���h��v�����=:��v�����������2@����a�o{�q9�Z�c�NI6�ۘ!��*t��y�2D�H�IEu���������}�w7Xi���m�9֙#Nɛ����k�k���4|ņ>~~��a r}	IYW�;:t�J;��p[]�<�g�� �jɰ�7o{�$l ��My;f��)X��Bdug�y�ъ����FuZ�|>�"�wu������_�zSU�yqn����F�#w/��;��@)��X26f�\��,����~��/ҋ���D|W(6�y�H�U#�f$\��������h�$�0'��^,N�s7I�Y��c����~Щ.'�7z��V �h�[\� C��������z���J�U����R�n�`�	ܘ��g���U��5#;�&4}q���zv�nr�*Y�-/;;�NE�������L��9�k����k/�WR9˿B��6�ex��l�p�� e���0A�6Ng�������0++k>Zf1�ĝ/�)zG޾~=.�Ń��]$�^'�z(P����lllܫ�گb`a�(��iQ�?s�e��<�M�.(B7߀J��O@�d�C�mmm'�ܖ�J�R�ͬ�%!!!�ďd
;'��&�2e��������談.��-��&�?d��>�!�_H??� T�Q<��c���I԰�#������(��dv���$حp��%�bv���k޲X���ݐ��n���b�YK|Ǟ�8c*9�b�%��Z����k�R�Q��tUN��D�����Rk�=����0ر[7�ӂر9azB�A^޹���G����|��bBS񔂿�lH��v O]{�W���a���ѣ""��U%�ssu*;?�
���*�Ͱ�����+ɫs�;&� -���H;�=�U�A��2M���q1 ϔ�(��@��<a�6�(- �B�y�8�'��:���~���c�y�2���rsk'iFQ͏��x�%:�Tm�G`)]����q͟���H���qU��5�N�\������c�`��f.Q�)^�����S�����ĺ@=��͛7����8�f���W�}����@����Pm$-5��&���2�7������C��7�S�t�3{T@ S�};`���"�f(w�{�D^���`!�
��, �ca� �CI��@V���t�d0rI/���#�\[H86�?Fߛ0��4��z� M���� ~G�PI�S�eZk��Ҝ��t]e�4;"Q��NB�#�t PY�8�e�'.���l � �!:,���Ŝ]��x0,�je��9gG[]!�)��7̆�D���<1�>M�:���U���S���PT�e��-�a��h�&��1�4�.>���k���a��Ҥ�֔Sa▫�������y��tk�Գы.,k�-7��ДJ����д5����{����ZZZt���TP,k
���g�e��^�[���:�*�1ekRw]M)4���5
>OVS��K
��/E���6��Q�WWh�����O��*?+�����ӫ%�߱�=��J4��~j�i�в�"Wd����g��VW�X�}2%�����a�H�I§�A�m��=Jf��S���?!�Ĳv�pI��Нs[�trn�d���G�Q�8�آ;�+��[��.cAj���������>����iu�~l+\�m�s�؂m�o�!����=���St/�8]9�6o��	#��Z�Q���R�A�k�����#ojb�$���H�Z4`W����s� r�%^�����҄���P0�m��q�3��u-��)��A���
.�8JGc]#���'��Jv�EpǇ��
@��~�ڂ�����������:��u\wcX@EG�rӘ3{{�}����m������uG
O�N���{����?s
۴iS�R>u�y�S�'�+��-�S̒��=_T�MO�qu�5P���!*�&<�*c7�$mB��u��������I����J�9�9(�5�������6̼{�N8q�	|�7Y`������eSɹ��:SIr�D9����~z��&�\{��&>�'��ݫ8�	|}�_fu^8��	Ұ����4����B8�0�����+ə�KI}̑�r�i�?'$�N�u��턂��M���ݻ�:Q &hm���]19K���Q������Kir\U�I{u�a�Y��b^�-on�SX4��&4E��Ll�bd`��	X�y���/
%@�Jr˥��&���$����H���t�c��#G�G.��?���kV=X�\�:V��If��^k���&�}<q��)I{zn.e�ȱ��P���z��%���s�^Qٓ��nJbl��Jt̋(-+�E�Z ��CJH+��J�� �1�ey89��@����gr����X��Ό[ 	'V�i+�)Ͷ�ӿ����k?1�)�J�b2�����a�i�0����vc1;f�O�y�]�ȑ�����c쇟{��q�2�o���HH��Οε��ov�ZB�'�N&���VV���c����ڂdD�I<��)MP<q@�Z�L�w�}q�������$������U��9g�LH��ٿ��*�g��tH�3�m�F<���m��ɓfR����/$I#���Qo�~��	7�Mtt�C�MI���{�#��~�:e�$'����03��Т�;{~BH-��;��C�8� ���=@�9)����j�[��XI����1,s�*��q9z�16v�G��4��ׯ/t9Q�*�;��L�X<A3S���]�"�wSu���ˀ�����"u��Z��Kz/ �)��a��>.K�%�����1	��+��å]Mf��s�Z�`�x�ǲ �E�W(~�Y�đ�)>�A����`bE�|A7�Ku�"9�s�z������sܲ+�#��=]u�Qz�
�஢-��σ�����2�t7�:`C�_o��^2�+�x�i�1%<�2�apf_ONG���R���\��Wߚ?0%=� .��f�M��4��w5:��x�_�c�6x�f�1��x���S�\V�y��~���+h?ߗ��͝ˣ����;�5�dC@ӱ[<\�����mN�C'�tS4�����,�Y�灌�����x(k�k�G'
70o`����4?�,�p���W�5��u�%+s�\P�|�F:v��GվY�UQ��XG�&�D���L�(~�9 UUU�5�������"�!��!�V��G�^JYk2���P�~#437W�ҢI�<��:��V�m���h�	�r��i�R�r�lJ�⛀-���(��L�
�h6�����t�$�dٚ��R��x��5i.-���w�U�	Љcs��������ǜ��r���\DB�hkh�p�v�ˋ��^B�`p��~!���O�<�Z��Ȼ���k�X��;UӒ���;���qT5I�;55�oe)��!h�x�{�:~���b�ƕ�f >$�R>/nb,�Р��=��9���������I��UWW�bò&g�n�Z\���_x��0L�3@��&V@QP2~6� C]c�sk�)�*�/�x�����`#x��@�狋��]G���oOK���L�Ԃ'smd\i[�t�}OOC�c��e�W�+�@��՞y���M�*2o�TvbH��B�ʍ��H�kbb"��S��N��q`q�~خq{� .t�JJJn��_��QMPXXQ+�	�R0p�U�i�iJ���1v��A���Ũ��>[,ύ�[AS;�O��7_�6h��X/��)ggY��ԢD � �6ܟ����� { ����z�5��^Q���������gG#���P����DRB��;���� �� 'l{�VOo�q��t!�cOu�Lf�P�]���$>�ܔ��S� ����ǴdZ���5�ʼT
�,g�>��d<�|��U|��F�7ǋx�e	�T �����4>��]���L�PRH�\X=����fDc���V�̑��߰u�	  �Nh�i;�Q.�Hv��'&îFZ8�9���1���o���<�N*�����o^�F[�h��Q{ "
rq}� ��	T�����&D��� 5??777�,��X�]h�lM35�"�n:����ԑY��ي�ˌ#S1�ed&&zz�5�j�2.<�����@�,"*�l�5����=
|髧D"����GB�(p� +<����A�]�_Y����J����(K�����ʱ9��݀X���E3CM	$d�T�[}q�H,r��kV�t�d�1�� �1�m��A�z0}�6���. T���`ު��@Iܿ��KSB�7�-�z@o�s��0J����x�wFo��4�v쿯"P��"Ö�T�9�������J�x�]�S���#;c���;��B�¼͚��UY��<�ݺmt�儦�� #��Y�H�~��H��Z1]W��96���@@� =>ell�d:P�$�-�,������.,���]v�f-��qph�,B�~������ܗ�s[��=1e�lk�~?Plˋ�f�i;4"=z�������19�p������.�qr2�owP,d˂�?}�x ��Z��iW�Քb�&�������)e�Ѿs��?��HS[��@@k�b��Fg���i[3�3(��D��kV/G����4��AفCPS,��F K�e�]��kpAEe����S�d������ �

2pu튧ؑ��p}�;/
�8�;2=Ҁ��`�F��,������̌|N�AHd$�V��Z|ǉ�<����S��@��'XM=oіb�P�����H�	$c)�. @4e�Fc��h��Ё���N��[�(A���5�B+�?��Ƣ^Q��R	��m ���
T�~��V&J��`-���=K NU��(��q&b���Q*��P���8~�/;��(H��'
j^��@!����dee���M�=L����� ��/ۚ���򠞖���w�ㄞ�D�A\균���VP���z�p P!y�?f�.�O $T�������t �xC+�#@6A���a �Y���/�RAP�����Fyq���U��p����/���i��;��V��on
3؇FB}s3ްQ/����ĝZ�9�G߯�2�u\�HK!��+&&fO�.��}�󡚗c�k�ݬc�E]�s=���L�5
���}'�g
o�H����iF�N��]�/�{���&���d�H��X
���¹���5D��u�s��=��d�Ri��"&������c�H��m���$Ӫ.��4Q�����;7w�K�|�hf캚��|��}�J���(��wbq��l��ć�#����kB��oV��r��dm8�Ҍ<�d+�S����}�j��,�S��v�A��D
.�𵷉��.%v�W���̟�`)�Ù�*�y���ˇ�KG��h�"9��ff��JN]����k%(��~US�ĺ��͍��8,��_�)�rVZn�6P��3��D�x��{h��ʌ��b��f,P�*2 ��ԑ��1R��V{KRˠ
��sߜE�"=%��PS�fjB���gED ���7r�f��="/=B���_�rPdi}�b�`e�w�6@ך�gI@ ���N��xT�cz|A�����)f���9З��&�$����J��:����(���(9�������	��G�Sk����V�
Or�Q]DL,��]�v0q���"���מ�)��a5�[�!^CN�6��\�h�[�`�&��5wEZ��*
W̧r�p%��D�4���<&�ne�p�@
h�$���:����%�ɫ�=c��jwlmǿ�b�@m1����^�@�`�	�^9hW�"�[ەF?�-��ʷ�w���Y�EY�p��o�X��^^��X��-ŉ�A�l���*lpp�wa(��|��ڞ��-�q�]@/�26Yss�:P���B��l�:���#�R�Q������H�]�����U
�A�����������N��I��L�St�w֢�sj�Rr'� ���4�.L���V���P�@������e�;	�i��&�SP"'�։/��F����*���s�Zbi�C����EN�Tҏ��sqm��O��ގ,[���P�)��:��8~���~���A^^��!�\��[��kM�&��:N"G�&a���]/�����BY��;�}e�ܕ=�t�Z�]�R�J��K��X䙮$�<��-�Vi5r����9��B""��Y��*/TQi��(�
��l;~(І4���]}�.�!@mp���dݜ]��z>PMO�A�B��u��e� �.n�=ٱQj�7��@(@�kR*q�ª�DF#�G�*EY,�����Tj4���$
�����7�UUrrl$�����W5�|i��
JX�U�v��Ya��P�,��Z�L�}iwK4�׈�4@PPPN+t�p�;��p�}��� (��-�=�ƃ���a��������%y������%1w��,��s����+�������w�?;�����
;�����U �[sE�+��}t����9�0�=ɬ�§%66�,L�A�WE����.H�i������V�Gw7P?�"���Π*nJ��%⮷A�C��{�V�HA�������#ᶸ�Z3���v﹐BD%~�ұ1sh]�K�E�;C8zh�C]8f�(�WPf�2-����?�2k��p6��H�V��FBA�S�p�?!!\��/3�-(�oy��D��qy�rbr���[ڌ�kVkbn���'/�Թt���)GtDP!�t@���2>ݑݱ��c�sK3�O_ZKr�M��m8�[m<U�2�$I�7��*]34��!�3�02=��ۏĔ�q=�4N�2�^�L�\�l�d4�˱>���"c�Ҋ��gQ6'�gj���;��o�ɋm�.�w�4��Kr��d��J����vP�s:KW\��$�"�lv7��ѕ�
W:^���m�I��r�}tFb�a�l�jՄZ�v`hu�X�� X��+��WG#��7����߯�Ү�����o9�)���c�ek�C؎��y�����J��G�7�+��O�>���8�فF����������5����k�_������5����k�_���t�V��]�������W�]�}��r�����AŇ�Q8�v�5(�ĭg�~a��f}�u��5W��Da+uh���ں��͋/�_��>n6(2���#;�\h⡮_�9��Ur�㫧�'�^��=�q];a],�S%�k��g�����9�7�@>��8 ��]��ø7J�.�W����T�/[�����Y[��M�bd[W�ye�v����������j��I���a�u�\?�A����+T�������-�����7EE"�$ʗ�޿O����ud�Z�����hLo v	��hj��tR8��=29��.�]mii�j�����C�_��re�2��������Wݷ�N�lg���������a���"˿={��]h��׿F �X�,������}��#�(���ݕsЕ��Jσ�ߜ�2��������xL�:���S��p�s,��ۊ��������B�$�L��vӘ���9d'7���~�:��]p%�+>`g+t��+,�=� ��n�֌�fp�BL1�d��N���s[\;Gq9iyy����<��K�_��w������.2a�5�p8Z�����C�J���>�E����2�+��ɜ!��f��׻˦)��c��W4��7�*�%��N�))^��0��u̘E~Ö���n\�~J/�^u��`�a�cBggmo�ܴ��� Gί�*>p�r��UH �ky�L��/�BNN���?{�b�����3�,�zt*�,�T�k7�2�4C#�IoP�}���+^���O�67xk���w�8�#�Yy
�=��K5<��F��XɄ�?/��Y���I�RUb3[>�����i�E6�O�91�}OG޷����l4�����x>�H�"u��y}a�g�":3g]�N|�K��T2߄�J�κ�4�ߴ�ٕ���S��IKh���(���	,���nl�+nҙz�19�Y��s��8Ih3��&�
�W�i}ZZw��`V��y~F
ɑK�lBgu���uO72`n��Ŵ�Lc�g��<u���Q����m3�I�$On����f�&Sư��[w�����qM��� ��6��gM��`�z�+�[c�q�z��q.uX�fWjv��:�~��%G�.�2�הQl>8�M���xÁ�t��QZ����7�s�ȑ
��?��E���Ǿ��1��w����IɑO`[�$��}�s��tU��N|Q��<��[G����!z����ZzzA
ѧ q(�2�^��I\���;���YI�9:?a��L�9m�ޯ��	l�z�[�#����a"��F��1�<��΍��.F?�庿�,�U>[YI���2}�٦^��h������yL����yi~�:"�@���r��(G�P��慂����YSϬ] sH8@H_�JO�^��ҹ��s�.��$�9T��|���$>P)���:�����s,.
'#G^���4ش1�$0�`%�k)��t
��	,���H�r,����G��1	@||}㫄�?Ǻ���Z�'��"��a0 ۀ�7k,�dH)�9rZ��{o�Ʉ�$V�I�.�jN�^��;B[�q���b՞��[����zN�9�r�թ޶�Ɂ�]f��L;�jC��UL��4v���K��uI��1��[$��\A_�3���UUU;�R�����Dyrg��f���ڂzB�z1��D����/�9���&����2Ñ�˓##Q�<�{�t�ˍM�ae��Q���_��+3���Z6��?�S܏�s���'N��%�	���YW���NA���3��W� �?������υB���� ӹ��K�f�K�B���K�W~��.�6
�2����X�A/�p���X�ڧ_�v�vt���\�_�ȟ���A�J�r�H9��³�@�9-d7 �Q��9��x�I�C;-s�����i��숯3(``�0�.��lRSw���`nq��n�A�_H��rp�����7?C���ٷڇ���� p��g�9��=j��{�.�k6��y����$8������eT^W�z���o|Sp� ����-Z�m�xWi@�� ��o�f��Z��r!��͝����c&�!�s�%/����T����\�h?`z��&&��" �b]�K�-K�Ƴ@�͎�u���ܯ|����\��5�=�`#��~��q.G�r=�2}z�8�x\-�	��Zd�'0s5����2쇴�`�sR���?���̸�j����%��H&�N3�lf bƫ��1
hn����Y�r�l�r#�J}<;���LbSh���o���'vTJ�"pRD�'��F�����z�	3�Ab|:r�1�� ��-Q���뉠�tTѽ�L�!X���~	��%��'џp1���z�L�#�����a����Y@�#�5\J$�w��yf�߳@�C�~� �+G� n��D���Jyz� �$m_��!�놑��#�/Dy�m���`��}�z�.u5Ӟ��xT/w�?��u!
�Q�H�)��(��dʠӘV�,|��,{|��5]sD�O�\�yǁ�87�l�?g.��g@�SD�^�ߌ�`囜}жn߶T�-�VF��_�o[
��W�x�F�~ߺ%lD�?NWq��ӧ.@�P�����i���*�D�,
״oL�;��HEo�Ah��I9��(��L�?�)���z�YK�藘�x6�5`d�V|�)��ǆ�77�D��^�k�՟n\��cP�ኚ]�y����v-�+���!Iʓ���o�����x���"\o׏����C���i�1����sg#d�N+|�`���ދ��X��E]n.��3��pc�����W��
��M��L�|'e�ʏ�z�`����??�A�4�;?=c���#[=Ж3�G��
)T���bTg�<�b�Ի��]oρ��b�o��%���q;���O"��C�����kʕ{��e%�>�q�"�=Ԑ5�����ȑ⿏H��zL��WluNĴ{iQ���G:�ѧ|��a��I����=Ͼ?���4�GSN
���kK[� �U�w�лø�m��ƌ�ڼ�L�ϴ��ˍP�N�Y�
'Ghc����&�V� �W �����><�����3� m�L~O���_ZG�A�s�G%��v 2.G-�9�ռ�>d0���."Ϊ~O3�]	�:u|ś7V3�p���%�����W��/	�p���G�����x� hɺ+��l�Ì�O��7=�_SRA��.s��@��.�*_ϏH����jȟ[hh�����W��4�(ޙ8]}3_���$�-�3��ҟ%j6��iq%(8�+!פ6V� 8�m)�
J�& 2�����Gg�Lk?.�Q����}p>B�g�;K���)䲝�AV����K�i���Fi�� oBBM�E�s	�Ϝ��Z�C��%~E2�I�2�3����{#�i����(�,�Z��`���K���@S����N|�w�<~�w!U��t���1#t��[�*�D���BY�?P�	SA ������v��u?h��} `פ�6
r#�R��W�5�w�o<��k;����#��x�	�jdrWMM`d�Κ���������Y�섓�;HuOxSO9k@�O�X�~�߲��3�'�-�z�V�����^��Ys��%�O`���Ty���B�/������'U��l���ɰ<�O�����b1V=�ձ^¦�};�"~������x1X�UE���
s�R��ݳ
g{���ao���_�]�qO��
J<���}��/�׊��b�]���ƈ�����\P���+���ֆR�G����*�L�GH|4w~���)����l�&<�Px�pa~�a=&O��ᬔ��_Qf������o=R�d���K�W��ll:�?��?�P�R0����&/�T�UȇԮ��r�p�:I	�ǒ�����G�@^n�v~F�����Q�b1�=�np���@-@^��hWO���W�S�M2���Sυ�{��%F��{� 9L��l];�|�FF�O�_^N�54"��8��;��t��]g��΍��")P����T�@e��dj�w��+,�@N�$]>,���Y�����ŋL��,X����T��o*�{ȋ?m�B�Vť�n�ޛR�N}x����x�:��DT���)B���B�OCA�
������j��yVz��"��*�\�͈;S�~��f��~��=m(���U��9�����Y��VX�#Q� 	S��4Д ��o�EF��>ߪP�6�YH)�K �1W����o�j�Ad��]�R������
]���b;�d�N��q�۷/�jzK�}�����!�e��t ��'m��0O��9�]�U�<������Jn��'���gCɸ�_f���]�Z���������ap�~!2|v)��]�y�N�S�@#�CM#�\ ������D%����鍛���k�p�]�e�<��S�q�o��pu��ug�-���#�}ߦ�uC|ӣ���GT:L��=�%�GhMw�3(.��.��q�^����6-]�@S��0C���8k�7��
ԩ���[0�؀n�g�Z�ᣆ�k���]tK�]��\��(��).o��n@�/B�/��-�k������<9�56�~(�<�4kn|�p�4��N�g��=>�~�eC�����鐫/���?i��Ht��y��4��jJb���pa�-T���Wz9��-r޶�T����
Bxa�S|���ʆՓ��)��Mk��e����v�W�
����Y�Q!J�p��l�:u��Gc��R����8�0�b����3&ك1���%�����G��TlvJrr�!;��D��bh(��6!���Y�!��t��)�y\����8����}�I��"��x�[�3�H�(d!Ş-�9�wVZ&XC�5�����U@�B�~@�?��}�9P�h3��x������#?� [��
��L��ߎ�V�:�A133;*&v��}��`�=���`�6�����*��7^M��i�� ��6m�����"C Ic4~�S��Y��m�cT"g�K���f��w?���c;-�3������ֶ�/AcٽU�ů}^��1/�< Ö���#@x��]�nN���@��m��fRo��� �[x�v�M��u%N� =1��%�-�s/�*�
	��5SF+y�c&e�L�p@�}u�E��I�g6N���.O#�I���B���֫���g M�Vp���v��JHL��#�)�+U���!<K�̌cF�!r�u�#��!�|������V��n�)���G�)N�V7�.�n�ph�dGnz:t��6��@��(-��!ZP�)(��G.ԱY#�g�V皟�:M,��X���(���^@G���)Zt���K��O�\�g-EU�0�~�F��o�����N��h�b/��U;Y)��q`��[�À���H �����<ʨ��!\�Y �z�S��$�Č_�v����H[�X-�u�����ɮ�8�����Ӎ����Q��)�X6xa������Mx��y�ʹ o��� '�1��� �'�q�{�۷������Zw�W��� *���桌� �ieB�W�1�����������|���.Ax����jR�,/鐀c#��V�����=�&聐��w�ѹ��_�ײH��$���6��G|u�@�o/u�G+@����445�	�o�
W�HR����q(w�O9k�Q�.��N�tr�:�_�&�m��"�2���Q��T���Nڑ������mRY�i)�R�eU�!�?��{�'�vP�u
���0�p`C^�&|52S���&&sՈ�NLN�m{V��"���۴n���0F1����Ce�x:x h�� ,�X�k	���ƠG��a��Z��u���V$�2�f
�@��u��F%�E���7@h{�����\ ����C�7�r	�A��u���q�@_'��u��a:u iQ9�<��D�7�U�ps��}�'&%}hldy�/ay��fnfv����@�7k�t�6R�{eʛU�E�H9��Ӣrv���ۭ��LL�X��rg�^����ϛ9<x����nn������y��ù�\\����ݣ�{~&�-w�t�Q����1�gT#���?�ʸ�Y 0FGG'��:e9T�2x	�ֶ��D"�꣤��Pci�adf6J
]i#�4��3pJ�133縭�.�,�c9��5W���g�#��U�_\g�U�O����=�\R��a�XaK������W�@�*p���94v0���(-����R	~�i'Gq5���L>�Q���Ρe͵���6^#!T�Ti��߷�_���t��`����-��X�G^��.�f�*��9�ʠqP�ޟ�����/`�[WKߘKɑC�^.^� 6�B#�<�E^#�al��26�������)�^m���MIz���:��l�ҙ��ӫ�o�r��@�z�$�J3�@�-���iyy�g]z�G��c~,V@TT����n3?��I�0CP�a��U�,�p���V=/�
͚��������E����\w����y7�c�͏�E$.�$��,.fK�,������<4%ۚ�̟.K5,���hR\�"g�W k�¥�E�s����o��ȳ�sr;v��EF��zc����a��C���ق���ccc���2�J�0?��%�A�����*�<t �G5�Fh�I�0+��b�Sh���½ui����LPPЍ[���behM7��Qomi�F��Jɇ^�:�0 r0e�
� ���yU":V��0�d}���4W��<x�Ӻz�	�N�)i+Ԥ(n0��o�j~����X��������Z�ڏ���o��~�2me����F͏Kf����a�_�C�F��]סC=z�&��ٿÄ�J��c7\]�����_?�m��"5e8����	@��+/xuqz�M���vM���IM�#Q���$�ι�n���[E����V��%��(�v�h�ў��͛%�ypL7������jj��߿O�	iYW�?�cR1��ۀٞ�w�e&m���k�U��)M�ἠ4��E�R��2ؠ.,3i	t2�#9�[���Gc���oW�LxXX�������|��\'����0�g7rY=���Ν_̒�s�n��*Հ���г
�D�ؤQ}�S�A�zyv��6���ZWns��
������7��U�^4��\�d{_�80=ҐC{9����*���3��#��q�ahq�*0DK���@�WG�����x��bF;�b��BH��[���9��!�)Cå��-�e�\���fDv�Ѩy!�`�#W�A/�I�Ku�H9J�h� g��"����,}�K+�#==d��	,<]���φt��eeeuƹ88d��������	�J���� �6���evc�"�y�9/��fO�Ƹ�%{n{���<s���@�{xxt�ق�j#���7��1�}�_�e;ԟ�����W�e�,��7L6<�}��5��w�LP!������}� �7T:� �<3�i�R.����K��,��л�Ns�yNs/Z���?<��}�m5W'��T�Nw��}[Hx5E�<����02�K��0��&��%������7�N�ŵ�gT��y@=������Fi��(yB��lMP��=���%��x�2�/�X�c�.���\�����8QC���"����p8���8�h$`�|�3odd��{F��2�:�ᨹS~�X�ŵ�������sտS���DުrJ�T{���"OƁ�����T�i��;+��(��P��9}Xq=�0�s�� �B��3�y�9�L�ʘO����S.{�U���w"�3s5��h�b�
�-�[��%U�ޤL��?-"�ռ����w�9M�>s���Qr���KK䌁�1�'k����E����@ wLB��:��ݼ�-�ե����>�A�V���,����s�#����/�K��O����W�5����� E=y�diQ~I+[ܱ�Ro��
Vʹ45�Ƥ0cq��̎ie�x���.u�Q�^��eC�u~����dB+���㲔�ᩩ��#v ^l��r�,��(�|g-P��^��`߾x2zn~S�}�Tzz}���) �R��,��w��\֩x�A��ȟ�8�*w���fzX��� f�������=���Z�n��o�FFge�t�~�<�~��<�~����D|�#P��8����U�}���q������x�@ >�M?��J%>h+2Y���I�מ���IP��G2��ڴ�L�'L��xM5%\X���m�l��~��@�t��q�����Vm�1WL
h�,gj��Z�~������,����.�<q}��NQ�yX��E�e�N�i��p̓	!Y|{iuha_U'M�K*{��?��N v�.�x��dx���l`r�r����5�J�K	N�3sę9������Z�����o��(���i��:�}�����lV������xu�.����WW����nw6�u��
kyw���ȋ�3�����9���!�c�����n�A��q=�c�h֜��:Lt�3���u����B��m�d��&����Q���a
�ؕ����B�_ЗX���c��G�Q�'��
y�XcwN
����1:����10�(�'�o��?U�S���n�Ҵe[��l��,��!��r�.���#S/G�_���r�<5���2?FĀ�x�k�4{[KGGp̻���'��x��|izN����L��a�|c�&U-��w���[���ńᖎ-IbV��=|6����R���?�K�����ĥ�s9��ͥ�.�6g��JKo��z�qx�O��ong
���jR{�%���7��E%hh�NGc0;�n�36�
�d4�����(�XT����ڝ��C�~}Ow�i|�J��i�W�T h�&KX����1M����]�⓫K�J�(��>$
���=�b�.5���m�h��TU]�!��U �F�Ek�X���@�z��`d���87h�F��8)����KV�[:��L�)p6|5?�33ުz^���z��S���#\��ShW�Z�u[Mw^�i�@a��l>�`��m��քQ�E�ED��D��A�E�"Ң��D�BQD�4% ]�*"ҥI/�#$QZ ����ww���ϻ���]�;sg�y����C[��ZP�,_>�����v՛8��l�?��1扠!��,�`�y�f�^b"�}b�п�okǺ!�R �A�P��>���*w.+G��(�o��d�q3��#N���RDb��7��Znl����1\�zL4������C�O��F��y�-���D�8e��˴�&�=Xw�Ծ�}&�߄�.Z+zΌ?6�<P%mnKS[[��?Eu�M����i��؅�]?�Jo!�I9:%lf�_�YXXj>�o���%�o�֒���Z�ϋ����/RR4Y�w��q�y�i3e��,(�w]JO�^�µ/vx��������P�����.��nJ�$\�����L���q!��$�I�E��� uu*_�И���J巬[���%zġv��=��뎹�s1'b�ί��7�zk�0��渂�()�K���{
{#@��d�T�L���'��s*�6|����Rn�(Z��ghCM@7���7���0#ed�f�CV�y���t
�_u�]��dg���=��6��]�D"�Q?>/��N��4�TC������x��I��K��w�Fb\��=���"�5�W����T��{]�
k���q���Y���AA�CC5Ք�=DT"��4/9 `�@�����8��oƾ/{o&��y�罽�5�~	��'��3! �>C?b�0�X��d{���X_�Cj�}�4�GȘ����wt�/�u܌rF�c.�eo�L&di2���3;�?=�������Mr1dM�o��{����R�"��aoMe�?m2����]����IIK�gzރR��O0
�����uuuE_b/r�ޟ��d�JZ��V�7��_����w�<=s,=�p�Q�� �i�^��W�[������'rʣCBB�ʂV�mjk��@5
��j�l|�Hq:���@]�|����w�@�s{�o��fW`՟@wK������3)[��u(�	R�~����5�x ���ة�f/��������n����.ԩ�䩳[�O���B�h�y��}���8�7�Ո(�y��
��>�J^��7ٿ�H��[ok�yñ�(�%\u�d ;!�ϑ7�;4��q>tֲ���X4�>���S@���=X��چ�6���	��~o�]��<��"��ѴγѵZ��"�4�����N+�׵C��%�U�▹��i�I9=
HL�>��j4�{�&<w�e�g ��/�	N�[�-Q!��R[[;�i�Ȋ����*6���-�n�j!��3�$`	����Z"��i_K�Ʌ��=K��V#DYC��?�-Ƭ�S��h��\�|*�N`�MrS�ZK��xW��z�������d��g���ݻT���֓�}����N ����{�S�}�]{{�G.o�2��ð!JK�0��_K&>��u�h����<�յ0�5&{}�hF����c��!/��|�	{τ�54P���F5p�o��i�5����
����}�����k	��h���p��9.� 3����oݯB˟*��u	;��
C_�	C�G�5<+,)_�(�4ɅԜ�Sn�;����r��֗z�Bɷz�\����&����5��vu��m3��W�&k���V܃.��Qc+��nuw�{��ژ���;���?:�vw�\�|iaq�1�"'f���zŮcw�d�C؋��~}A(
M%��\��)*�}Vqđ��k������v:�GH���鱎�wCI��&υp�!|5c��e��ݝ2������`���	(�[�neQ�$��R�;U�?� j>OS��O��R������B��,���iu����|S��(��V������$(G���)�f���Gȧ$G%J��Xo��!4҂3,rj��(k� Vu���U]|�3�"�t,==��|ԁ�3A]y�JR���-o����k���O�=���l��`���d�TB�]m���3h'�Q�eC�k6�n���I�NC�O�%0=P�X'�S�e����7�$d!�cX8m�d����W����0K�h]��@�BM
������z�Р��'|�����VI��xܳ�l����8c�V����7�h��^��7����u�����'=��gM��Հx/43�a��܂=�Z�r��S�.]���I�佀��{���Î#�l����������r,Vr�����g��6�zLiR��kǶ!<�F��,� ,[]���7Ht%�F{��x��
!�u*��٭lG�T��R�v�}�-sf��&qB�3��j�{�B����!Ή
 X�s&ȑ�������w`�1����ӂ�-V�yJ��w����c�� K���!L�J3�i�u������~��N��������0�F��H�5����VL�~�Z_@�\�{K\����ys~7l\���0�t��8X�u��2���xgGd�*�Q��(�5�{1�e��p %j^��)?)��vloԭ�!!��éAA�P^��lS��aS{���yB�8H>wNd�- �w��m1�d]�迲�R���~qI�^aT݈��w%Ap�2栂BZ��݄�� �~���Gf���?==�7��E��
��tS>6^_��D{u�٭�J�%e�pq<�q�݆��Zttj��t�V���鱧O�N5Rp��As��[�8�r�
;`�gZWw{������`����
����G�n�����g:�3N�n~�^ P������|�VX���ި���^ D������] ����N�o����%�-���6�{a'iill�'4��Q̋1�.Jyс��;�L�:h��{�Dݤئ��B֤�fᗳ|
q��p~��X��\�������\tr�;r[B�Tm/^ԃ���P39�(^�����]��2C�h�e5/�s��͛u��߯�L�FVC�	L#�\�r"$���gS?D��zoE���^��e6��Q��ܜ$ e�O@�1�I,cvX�Q��@����>�����Ȥ��PU\�3["֣�e��o��B�|�����D���_r��<��@D�ګ�.��1(�
�
������A�bM���[Hǀ<��4J/����y��z���n�Q�i�1o'yܧ��5�َ�4�V!ڟ�	w�>��
!ni��>b��Coj�7�K��+���ͺF��$-��� @�
��LZ�E�I�\�z}j(�D�����ɜz�}y�稙�ݕ����yo:�m�����q��z�#��22b#����qM/;���`���yiժ���x���kFjcF�
. :�d�ZS�/{###Y�Ik�o2������LяE�{�!��#(����������qU꘵�Â�T᧹�ƊŎ���X���|�t��i�%�߇{gKbۏ|�ؤǊ-G�	Y����z�a��N��k`�u�LMM#��L�����i���bШ��?�D���`�G�h�b����Ks�.S6p�g����_WW7�LKNƐ�P53}������i	F�[���.픐�:J;��t>P.�A"��7�\�����`�w�n@B�[Ն����PH�0;" `*��g%��GO)����~F|���s�ﺺ�5�����s	0t����.]x����@��`�	�c��H�3��̸!k�V��u��~�m>�G:5R�����8_��[ҽ~iߎ���_��5 ���̓4&�w1v�T<_�_g��]8=�B_\u�f+� Y�:U'M��P3)��j�\����dSUk A��i�hu@�����s}�,�����<�9LJ$f:]�	�	`WG{KvZz}�_�,��[�K����
�opT�8ߨl�:�H}��=�|�C�9۶n���ܣN�b��D0Ӿ����u�S�!`�jTe���f�}&��o��#�����8�C�� q��q����7��!���ٗ�
|{f�!���9������������5��Fs�s@�؛g����.K��4(W]&�Itvu�GH+*��Gu�j�F��H�~��$�+H=���~hW�h��鐛�������{���H�al9�ƥC���`�Ϝ���P�ǋIқ�;�;�_����Ξ�
\*��u�g�jC_�ټ��/���������]�1����=�����|3��+��5u��^�)�nin�4����Ä�Əz�ay���]޿����h����{�����,��o߾)F?���_��6c�N>?U	��ҍ��?]�k*���U�����\�Gk���,��OUB>������GrÔ�_U��K��
�B�g��fY]%컟Z�pl
�+0��2P�{-8F,|�Ǖ �3�ж�܁�%�yw�^rt�r�wS�
T]<�4aY���U�.}�ζ������By��e C�+E�+���ۆ��*u�����?������ ��{�_B"���:쒆2�y��s�g�B�o�#��>��-�4�.�*��� 6��d$b|�p cr����VUU���ʪ��vx�@���Xk�\���Z�[h�]2���V-JG������ �8�'~|���C=)���5�����s4��%fA��I��e��Y݅j��3�[����b`���*��p��{�F`�q\�Y�؋��?������ŷ��=65%���3���Z�e#����o��0�܂��ű)��PVi҄���W���V�'�8�#�y�;����xR{��(��LFy���.Hl)�s�u�Q]�P}CD�����]�v��x���P�|�A���$+U�U&	�9J�ٝ���
Z�雕>��"�����p�����W����$|c��3��.`?���ߏ�e�F�4Y)�nj����)���.��8����Ѳ�	eth���5�W�Smv,���΅b|�|*�y� �Nd.$�81�jgn�X�����k��X�E��!Y/j�,n}JJSE��F�#�Ҍ�AyHe��-WG�xs�6��A�L�$f�;��XH�SH��/l�x���Ok����)�G�oL�MY�&�v��GO�/��1���ooqDW�K�_}c����aA�Lkvl^{���Be�,����D!�U1��d��M���U�%z�L?5��T�;_�����V�v�Lo��n�{�';l\�D
j��M*&�V�<�D B\.W(_X�MҵLFRK[h��y�ܛ�>q�sd��v��Ou�����[rKOc�dt�jn�B��۟�<�)�k���|M�������)�����؄:J=d���9I�g�[&����W�b:��ú�2��Ѕ��Õ���a];_�$���C�kWb��+�OsRx{
�w~�^�����5�k�v�op�fD0�	�t^�:7Ӱ?B,	0�[�G� �I���M�+0P?}TK3J2�W��X�`Ҳ=p� �P��SY���JY��e�s�u	�(E��Q���O$�,	"#�'K�É�L��r���x�|��Q���!RA�����pxY�ly�*DX(��1=�����zƈh*F�^P�9b��p�1r'ށ�������T�l		�q<F���6r#�úLV�����1�%�cD 񔯻�O� ����f;[��}�?�^�X�Jr��b���/3���ZЛc���7hu�ܵ�����&(k3U�������_)A�-��C"�g����]��3���;�A@����a�)��g�f��ˢO�X��48�v D����ta���L�;���_C��^��9���u�p����+��Ϊ�-7C�w@b�╏�e��1m���Z��b����)�xns�z���y�b����Z9��}����mY�#����)��1�ř+�*0���7����<m�����.<N��ZYT	��FҙF�hj��(�|ܑq�(��Xz_��@ZВ��.-ŵԻ���Z%�H
؀��Ɖs\#l�3��w�J,'�kS� wf������q��1��f��;�{Ӛ�T���T��{��}��94�I����ߓϴt=׋Oc��?�um�9���
�ak7�V����9�K��U��<���)�x:i&]�x�ݣ3C��I-�YmS�k~GՋD�g_{�֚�	N*3;`���J�?F�Ҩ�ԵX�o.9w�]j6�`Պ����{�ˁ��1����u�e4�c��9	����cF@��w����އ��q(�L46�%����9De��ghX2��$��ˁ�����-/��pYΫ�[�^ڼu����]��v4AI��:Z��4�H�IN����������SY�fs�f+��7x��&&M<&4t۠���FJ�L���f)�f��MD�˷XH���r/3I�_����'i��[o/Ҹ����S���X� i�5^��1�\\���<�߯����ŞH�TA��X9�� �L�d"�l6���`�׺l��[�ML�
�\���-[X�u�x�����aV�m�������� ��=��ܤ�)���M�'R�>z��P���}����Lʦ�f��*ڥ�2�d�G����e�Cw���d9�y_����0Z���\�Y�G�����j��V!%I�)��h�E�H�p��ǟ��/<^w�EoAkB��L����p�B��j6�`R��H�X��:+f�ivs�/�џa�5ȗ��� �Z���x�1���D�?�S`j�D��B�,�������4~]U�F�Ի�Ğ��d���5w;$$��2�T!t>P���~�z�+��@��)*��௣D�b
���b�ⶉV!S��^)�/<f���e�u�3fC���/̷j���;h�=�j����i�{��{�@�x0v�uo_��kCGY�Jڛ����7��+'��`���J�����GT�j$.q�����'`������(O�ӏ�䄀l4�Z&�]�FN��/_��U�GM9d��x�^}:����iuX���Dr	�4"\J_-B]v���V[)j��$�n���� �ͣ���Ew��s����NH��?�¾;�$~)�b&e=ºl��\hP����)�sױq�Mh|�� l���<��)~.�7۽��{�\���I=sQ�KS�.c��:�=J��֖o�]��E��9��K�&�_�P
_�۩����:��iP���x��+]�S׀G�r��{\c�n�r%��U&�y�؍Uխt�iVK��_Ny�bXQ럯�W&%`}�[��6�'���H�;d�����m4�҂�R�����Ǖ�2�{�{��o�4�A�Ŷ�簮d��b�lt}�vѮ<;�4��*��̃k�f.S�����$����e\�Ju�]�U��2��/�Nmu�����)s���S�eX��I�ZD�u�]� ,fv�=�}�[P=�N��?��`�� ��q(uj�%�BEk^�\Q_W7�Z��n�i��j��s�W��I	4��/3�[7� hֲB����r��P�.#��`_<�Ӧ)��-��.c���;�M�7�J��L�{�w�����"�;e�o� ��m��8�K��j�a]}���Y�]B ��7��Ն&��Tf��EA�MG�tc(T5��������f�X{h@�z��~��lZCsّ>=�d����_�:����S�8�N�+I�1*���-̮�z~�����p��d����ӧ�H�U����^�n�Iޘk)��R� �^���Y�.HP��++K7vI
������w���L���<s�P��f�V%~�vXW�_�Y���ѽgL%[ ���b	z�B���O�Ի��~4}�c��[l��ɾc�����~�>�	c�S�S*�Z�O3T;��!�V�<��ѣ��Z�A�Ԏx�� xR��/l���HfP3�.r�z�d�/]E�)T�OP��5z��I���?��أ4�f�F7*+����B2vF�UG�tn�x_.�}\����1{�<~+|a1��g{х�0�_�N����~V��U�N�VU5p��JzL�Lyo�ݓ���{�BX����[t�n�ێ���#/���Q�҇�п(��k��q<�/r<W�)�]x�P�V,x������3by!�ǭ4.�_����r+b7+1�AE �h-���r����u�]�F8�<�����$k���Y	⡠�LGEB�����;>�A/,=۠��ϰxC~�O�׍��i�`-�P3l�՜~a�h���3p�70h��[{\Oﮖ���v�Va��/�.�}:բ��^3�	"�q�I�M+fP�f]�Y@��_p�K�Ţ�?�f1Oܤ"V!:���'�9U���@�M�h��� 5Ж�&{C�_�zl˟l뚾�W�V?S�;"Ϙ;��(��'xȺ��(<s�0v�^�#2Uqv��}b�:�%��/�޵Րy���y����L蛕455Q�
���ь��]Y�9�3����ێ<�ΩC��v<��X����x��YK *~6��.J������9�cjhfߙ
�l!6L�eW�
��6B�pIkd�V*#P��Mqȯћ�����-q�K8����M������8߻4�fYaZ�\rN
qWN���o/�ȳ�����*	���b]��O��$�Qܶ id�*@=��@T��[�V^g*���4���t'u(���M�Xp/%3��Ų��)�,ـ^�"?X�$X`��X<�OH=�؄P Hc�ؔ��^�����w�{%Bǀ�+�G�Z4�b�#�=�Z�3UΛ���&�]k�o�x��FP�Yd*s��x��R#�m�dd$G���?���=�l3�ʟ�q4G ��=��Ͷ��$.��(+�j�#�<�!W���:����D�����K���.�l~������hI�4�,�Mm�'�4a�aR:�sY�''Q���?���2e�����ȓ�8��b�J��Ӥ�c(یn��4����>�Y�M��K��e"�Y9e������X]������&���V�Ȯ�q�d�����]�v��(��W�q��F3�'����H� w��M�ꒃ�t����W�Х]�%��������!.��:��K͎�ʭoI>o)$R����e�3�F�xB����>ӵ4�u	U�ka7A��C=��4QCP��������%3��_����f��p\��Mɲ�s�G�Cf�W#�u;�ު�������V��cO��0�R������������[����~L�3U���z������r"����w�+1�;Y�C��c�}�ԹI��ʒ��85�X9�Z�j��V�]����̆T��jra�>��9j�������>�*�_v_��z\(�tڜ�g�8JVV#22Ȓ=�I|�	̏<�i�)�ׅ������*��ܟZ�ހ��D�����I��N��5u�n�]3o<�~Hj�[�G"O&x��Ҳ����,nwjgx����v4�����;�l���P��-��1�uc�Q��O��,�s��O��JR���d6Ӹ�LpM�u����wcםH{��S�]�"Rw�G��Ξ��0?]_/�d�z�xb����v��B$����.����m5�W*P?ch����@�8��ľ�{&*ǫ�&�b�*���>At��w���>�T��=��o6{'Mt7!N�G��^<��d��}'�����������$6�&.�����4��ϠK�I�;]��y�����lX�D ��g�s>���b�-���Z�
M���ƥ�4�����A4�ps\� ��"r��9���/Fe~Q��{-�u�\��d:pZa���zj[����1k�-/�+Q}�Κ^�ͣ����|�<+�1Sf�k�k�@��$ D��ѳ�t~��uNL�G�/NqR$)H�Ɇ-�|��+nZ�@��x{�6��W����g���`�V�;���z�N���;�����Lk�o�J
�dL!2�c��0f��,~�����U�����9��^I [��mJ6y��i��`�x�I�J�b�/�{��p�86a]}�5V_C"4l�Z�%.�-|�2��O�����M�Da�z��I�� 0Οyo�F����g��=�*���G_{sf��EC�G;���cd[���!�t!�h	[�ߤ*l�C��2U��{#��fU#Ǜ��E�����A\�9�b'�������Nd(j�����Br{�y����ĥI;��Qzu˗�N��)w h혞������ˇ���PuI�u����ڕ���D4��h'�pCp6+� ��=�+���!��4O��	�%@$
�Q����OH�_u� �_��r�#����]]]���(%����ݯ̱�?�$���ؿ�F�5�@0|*��:9(ɫ$%G��b�7ML��]�@lʥ�p1�D��+�k�I�>3��}�Kr

c��Uw���h$�V�/W���Z�uu�ۏctt���;�1xn#��P\�Q����fj�_<V�!�'�E�&{`V˂�Y+\=��U8��})�:���L���#�����SyGy�X��3�	�c�	y���iх1_*^���  ���mk�]��y$2��b�c<)�K�J8�n��q�kÏ��+Ъ�� wL�H��Z-�T���u��:<��8���͎��>���5��=� P+��0��{"�.h�,`1ľR��e�{~�"��E���tH�
����tll��PŞ�پ����O�\Rgn��4�F}���x�=�2Up�*]X;�:#�d�f#��_��DUo�dz���9R1zL?.1�h�O|%�w$�k� 4�U{Kh�hm4� O±�s�~�Ɍ"�����" P��v����
D��r����u6�ɱe�*�������H��XA��-�7��3�yOA��Xd��Nd�X1�ú�F�G�.�O��)b��<cJ���}C�VJJ
�+��%���u'�4�0_S�`����������e�
>�mZIٺ+)����� >ߨ�c��XP^�ق�u[ZZभ����,��9�}���[����O��Ɗ��ъ�l�η����#����SY��@��v�6���n�[<1�ݓ�-�Uh������>��X�rޓ'j\\\���n�(����1+Hv�}R�=�}��-�@�#B%a���`�n�O���ā�ٽo��<��S�Ͻ�]!w�V�mUp�a��7��<��C�h� D�ӏ���4qR�Cr�+�|޳J`�4`�������ɿ��l��
8m�G��]���g���k�M�zDw7W�T���s��]�����P`�j/�(OLq0h�$��"�S�І����	����w����"`֒��N�˞���~h��z{{�6���B/#Ș��[W�����F��׾�i;�-�gl�'�	�	}��Z&�ck�5�=unУ�Dn���C���'V�^_��5
�e���w"Os�!�zG�"��/h'
~gx7��W�����/��G�Ȉ��6�<ȹ�ZU���w Dp�����C&�+�	^W��;\ I�:��M���q�jd����{�A�K�Rp��1�a��� K�9��U��b�?/�|z��[x��Y��T5��v��ꥡ�>��|ժ̘��H[�M���9r�'Q?�T6`?��������/*��D����%�iR�m�zW�~�K������b���2Vi<��w��]�����c����Ù��-���긨�3����{~��4���D��cu�z. -Ȁ��������=^;?HeL�1��5�,]��/P�ѿ,�I���~��i5����8�!���Vf���rQ�s��e 7R�xU�.�,���M��/_^�� ���X7Ӛ�j�IG��z��bJ�[GA���L6l������R��vI��0����t7���ޞ�[ ey�P����C�7ޯ��/q,���[�����J��@���� ��s_�?!@�#u�g�ܶkè��4�.O��94 �O��Z3�Xq*KK;"u��H�����k8)��ǲ�L�{��W�uv�Ȅ�a�^l?yv���,K��mPPtt�}�cs`��o���l�H���0 *&CSH�>O6�!y;�������cFH+��7]'M}ֳW�6ڤ��6S��7#��mcG�&�Llʊz�p�`�i@��=��q+;���y�pFĚ���T���2��ߺ���já���U��W��8��_�����_@��ϐ��CV�<�䷶�mh��I�m��3�cʁ�C�����s�v-,&{خ�����{��,�p�"��������u�O���t��x����U�}��
e�B��]K:/6?6'$��b��W{�0��]�e����CGQ-�PEv�S����0\��k�-�
�z٧j��oι�D4 ���U �1i�/P% ܕ>�en;�-�@<�Q�����,��L �;�o~v��4!�VM��K\�h���<�Y�#9�����x{CQ��Ccw��t}�-k�%���gַ(�/	��#=,g��ќ����p�e���������c�3���e��_�Yy���*i�ߵ���yz#�4��a�lOj"�o_���Z+�A�׋}��;`��ĵ�M�F��М'[G�O"7H>ǉ+����.���Xc�4o�ܕP�UX�.#�N��Ӷ����ٵ�G�&,�����g<{o򝛟w���ԑ�u�\}�h��d�����E�]��ώ���r��ts<۲�?d��5���1�@+��n�����|LD���;�,ML�H��w��"��z`
���'F��j�����7 ��J	�Y�x��E��>�5G�� ��p���c�"�p��7~��υ�})���t~��'V��w�����Vߜ�,�g<�u���O��^G9#놮�����<�����ŐU����)9f'�ǃ��ܱcٍ�^�<�V+Q�vj�k��S��-�v��ٵ*�����8!�h{���aQ�
��ff����.ǒJ�l�*XQ2}v<G���������P��!����oTp"�����>7F��� ���?���6���M"��F�v^4��N�N��#)���Ti6ǗH3����ի��,��/v������jq;�6�l���=���oe<�@�`�}�p������&��GQS��\/�a?�f�]�aߙ���پ��7��\y�i��&\�x�x���󨍯3^�8[�f���6�K�]�N	�HhaY��y��+��Rr��#�frl����i����ٰٻ��Wꁲ�<�｢�ٰ�����j}���M+���$�a*���km��[����ǃDt����s{P�-�^I�??�)�z472��,>�w(#	�<�˰�kQ/6nJ����G���755%ќ@�c.�Z���1���[�f(��-Q���~V��������g�Zt�:xJ��� a|��o�L�]�3M��������k%�+��_�Y��ŠcEU���$܄s��#6:�E�Հ1fl?R��
��/�iZ�U&��B����c"�B������%�P�W;$UA�w���o�=��<o�Q455M>��~d���r٥d�	����b���Un23<I�jr��
:i���{f�m׿Ԭabڐ=�IK����`�����x�裡���	^~����b�1q1NS���P�􇯛��:]��8WĞ�������ѝ�]\�95���C@�]h�HG�X~~��']`J�>��!g�d�
�^�o	l"�J��<�{C�~؆�y���C[!뜞(g^�m�Z[�P�uuukAh�2�i��]����1�qɇߒ�V\O
l����0�a[=i��ȝy�8�ݚߺ�o�E��f��{ݛ�l꣏@�8����_Ȱ�6�A��#G�<��[�t����owƘ�;yԞ(��<A`���B�z�
Y�UDv�n��+�ڛl������/ @�(Sp����_����|�Nf�"���y%�}5�	f%S5�ZҏkP��}U����D5�o}�?ۜ���I���rv�w|��+�~���e�����;��C�X?�~�����}�`K�ݺ/��xU�e�q�9���5Chu,ܣ�a.t͋���?�5X�@���&�<ř}&/ ===��5��ژ�Z��Q�1���=G�9�d�ЄlU�.(lC7�q����w~��$��JY|�τz���?U�6�׶��1����ɡ�hwш�����R���IN��������^=G�&�B{;2"��Q�N_�Iܴ�Z�Dd�V*�U�݌�;-m'��@��0q�F*���B�oZ�^b���TP ki*<�mkk�	��������C���7���r�|�[f/��p�t�2&X���2�_���#�➏���oz`�/��;�:p�B9�{3�5a�QBB�0��Ө�kkk֚�H��������5��F�o� ��%�|5^� �i� N�Z���{�s$�-� �S�f�2qf���'"}�uԡ���݅N�D�%P���4�ı�����E�/J	��
���a�f�����Y,��eYK�/��Z��+��m���6���#�qd'_䥾�8�6{Ay� ����#cϾ���>��,��<�� ���.��R˔���6-@��x���%.�'2��U������<+$�<s�G��-1hp����0�o�JN�X��:E��{P��)��B v�E��]��_��Er���@�}�>����(��ܪ�JK=��EG|��w���5��S�(���1]ḋ�g����ZX�Lᇩ�%�CBC[`Ж�s���m8�b�c�^�$m�d��=3,��a���M�hp�x5��� G;�@��W����Ad��o%c2Oe5�ys�$�O��U���)-�B�T؀�55ZiFI������[���u�X�ӱ��#�6@|�+��v���.���O???\��c턵9X�o�׈���Pg���*��1~�����������'s��;a���]ԃ��V>�@�6zl~x��.n�Y�j�N��`Cg%��u6�v<ƞً����N*����R��|�Y�%P��)���Gy��J�p,�t�d�Y�b��;��w���E���iG��j3].�_�L��^����;�c���������T<8����*P�����Ϩz�'��2��k�����)((�E��P��-���� ��R�����]�v翇|�8(���QfK�y��v=���֬=/��5���t&���!���%�"�\�HFK�
n��"��Z{�֭�]&��t�x����s��n-�����DOy<��ÍR<�=B�)���y�]Ŵ�iW�|�m������>}-��5��w�	�Қ�j������>�^���n�v�[@����O4���|�1����� ���yƇ�SB�KG$�+�ץ�?�QO���ruȚS�@p��^���K��4=���@.���Ju��F\*�=bbᱳ׽�\��6i�;���ŕ�O���K*.V�w�CH���q�����1�Vd4��p���z�����z ����W������:&V������\�$�Q����޾y�r��!��K�=)���햾*KK�L���܊7T�^�պ2w�� ��l}܀LA(��z �"���יzT��Ɩ�����15i S�P�q�oie4:�;m$�����rxs����l�4 �5�\A�j���+��әz�� �����/~�>�**hD��ԅ��/��n�R�m�
��R	�V��Z'N�MJ�i}�EN;i2�1�R���6���S1�g�9#ss�agE�莤n��*ǎabq�	\�3� I�Мy8^��9����~�}��.u�+6zp/u�/m�~�e����Q�`�q&C��4Diy~�uW���"��"Se�[�' �N@��M`�o{S����9�I �����|�'p���x�@� �R2.��+�f�L�B�UP���g2H����Kv�"k!��a~�!�N7� ��D��.8
��NZ��4s��X�(q���e���ڊ���R@n_/X�}B�����tb� s���"�4����J��iR��׾vtAt%�W��R���G�]�f� k.����ȓ3u!�.���3�8)�I���8k&���3���&�&�j.�����t��b^�Ҙvř�;ԲNe?mh�\<���� �/g��s���zq܈K.�*#�5�:�knG�4�EǼ�ĉ�ƘO�:|!X��6��8�I��2��O1dSO���NΕ�}�ht��e���9����}"���w�H�jj}gG�C�{�\�#-�������c�P~'�fCy���`hhV�Y�^m ��q��db�h����!��~���Z�|~��/@nX�5�&�������q���q�t�avd�Iځ~#��ct�N�+�2\�ӿ���'��Yq�b_d�v5�Wq��/�:w��o	��{Rb���cpM�F��T<=S}�8↸mt�WR����Ne��p��������V	����%�S�|>ϼ��Q$�����R�W���g�L{��׷���{��N��x`^s ��ì�Y��������o�����@��?.�B�`�u����K���A���&�Q^Cr[�	��A�9\F�sת����o��s�a���}~��ܴjf,�y��w��;�#n�B�s�@�m���AF���w�f9���d̄8y]�x��6	�z���d9����.��U�`���RV��+�ȵ�N�/
�Į�����{+,�ƇX�r�J���3��f��Dva�:�5��<"�5�^� 	I�~�6���e}
��%%��+���h$d��|~}�.&��<̋��P�8���y]v\n�sN�ͷ���YD;b���Q��Ԕ�9F�J�KɁ�1e�E{�G^-z�փ�T��W�$s�M6H�c#������+������jv�ڎ�?CT�pX|s����bDYzW1�����#��PŖC;�ġt�w���s:�O��T��@Q�'2�3�:*�$�Tr^�R����Y�;u�-]i�!�qX��1��`goJ^�Cˮ	�CI/����K%�3���@�˴��s�`�A ���4_��~������B�Hԇ�$��H�����ܖu�sy��a�Z�ܧ�}CiM�VVWAt¿X�})llp��Dm���UYڜ�y�M��^���ALI��m�o����|]ï�R1H33I�k8�X�.N���E�iP@�p�������>�F�L�h��@̓pl{�;hafR�����X�8Ż6(� �x\��	g��ﴅ�{���nˎ��6���>�l`x�So��9<2�}�BjkIӎ�s
��ɽ?��3�]GGl^�O�U�<�j���{I/-��f`�|��a1��͍Z��!	����mY��S�{��������
HVq>�+����k�S.�2�_����;�9���
�@�L�d$��9Ob�Ĳ<���l*y{���=ޏ�L�(�Fhx��{g���[�)<�a���ʱ孒7�i�@O�
*��	������z���e��@�T�p� <��+�����DJ������t������y�Ӷ��Zl|��)����c_�1�9�d�Zm~\�˗:H�]���a&��PT.�R��F�;�.:�������(6F�{�ܣ�Uxe�����e��f����v>�b�s'}�d&Y�VA��̡��;P;�@j}}��u	�a�O�`�����+3R�[�1��;,��'���,Oک�ۯq��(��6�a"�&2̔�v�c�n̉i��t��2�>]��"5��y�Z��?�~P���(��P��/!���qH���"(�.z�@_��]j�x��^�,ϊ1$��`�͋��W��:K=d�_���J�^���>��WR|ۗ/WHHJ����+4�G|,%(���~��_��h���-Sߕڑ�·E�~-��ƪtAm��L�Fog!�d�Iut�;6�H������X�̭�?��>����qڕ������z\[�=���!��ܢo'�_�_t����u<޵~xC3ܧ/��A��\����@,�&sk)k��ղLr0]��$��ԹE��.�~�C>�#+�^��=*7���9��s�y|��@ˑ���i0���MMMp�q
�j�c�\)�s��d��̓{݆ÏJ��:��Dq+���[������|����h$�p��x~�����/�\��}�5�Z�� ���]�#/�����UO2\��NŜ9���Ͱ�����2�@;���۸�� Ptq}���8�������=��VQ��N{�ih7��w��C]%��.��]�XPx��م�7��&�#��#�:�j�#6�Vw��ﹾ)��!��BZf�զ�cZ�=Y��(D�EW�5G��ޭ���M�5�S���3*xT��.��h����++T�ҁj���>��<8(������������}�O����*Y| 6�D�j���/4��:�/���ºz߻`<������5�.a ���-��@%*H���*����f<�O����S�Cf'�[�
j��,�Z'��jx��/q^j{�<T	������)�WǇzt��~�ւ�l^^bd�f���%�T�o�d=�?�}y<�����h���JhWYn�i,�-�T*q+�B)c�$�B��d�m!�$�J���k%&��31���y�5��=��ǽ�Z�9����|��sX$��楻\�d�k@��*�r�w�u#�ʜ<%��]���ӱv�|��J����[Y���=�~����,�,q�%�5�ǭm���+�:���[Y�{��4��2�b��\�/�.i�Ԃ3�ks;�*���N�Ӕ"�O��?�C��\���_i쑸�����S�l���<�H{b�ܭ18�������g�z;1��3 ��ܳg�_Z��������s+�c��!�3ǭ��
55�� ���Dj�hCѺ)�leᵠ�~��u�wÆ�RU.d�S��	�͛5{v���C�2��<*U�����N�z�KR�e�Mˆ���S���C��h�b;,�p��o�Ǿ-,,�������Z��1�M�[���~U�ϳ\=$�96�%Ǧڰ�g��z�?�����~�˵����1*#P�Gc�l��+ѩ�D��K��Z�q��h�`Og�����tK܋�'�l����K���R �IiɎt�p�I��L�5�J��!{���v,l��Xs/�^�N{�/�I�����#�1��Х&�?��9�wL��Z�t�KC�?u��I?+�T�� k��7D/ְ{ᡤ`���F�O�S�V�� �Oi��K���)f�譇x�x��L�h�{�k�%�)Ē T(	њDe�_$�ȉ{-V~�w�$=߂rF�Pe:
5]�{/��s����by�6��,�iגy�,���P�I`�_rQh�L3./e�Z�gm���L�q:'W�&��ʝ�;m���h��&u �����Ց�6l���x�Q{&��L���6������nbϟ??WH��]��~׸���x=��h|{�	o��O)��iO�p�Z�}�@�K��90s%�Q�/#B͑�U2���"���Y%�0QM�~qz�\�ZL$�{�K�^]�xɆ���^3�zj�.~��egž�}3�[z����Wo�����)?����}�Xí���S�;��d�v �m��`؀��fe��Gj��ok���k�8�U�y.�E�W���N��D��f�)��R�mW�䎵Y\F{Fx_X�����q�U�*Io��¸	2�6��~^�ô<8��(Ԧ��?�dտz��>�Kպ�����ə��BK��m\<b��_&��h���_��X�/2�h���F�Q����_�gDd �)]�@_�'�i�S��o�����ٽsa�������w&��۹�@�/쪰e��d��>�,LZ
����:��qeG>�~��൒��d��9-��!����#���ܣG��Hg�j���GqMP��3����#�m��}4���F��V���a����v�ٮ�B�q3�2���q��(�z������$;a[ҋ�qn)KQYr����=��zLS8)���l
�b�A�y~;,�B?��6i	��-�mS/a;'Ñz}�9����X(���=��u�P��͠{ ����G�]1�;�$-Q+sP�O��I΢"w![�9�b���bEXV҅��@y����.�J.0�O��ߒ�]W=�gI
o,j���;z S5�x?w��9ڒ��'�a��i=0o�4r����Ց�������M���5�D��^���Q�M��t��^
�]W�Y2C�wz��WU#�' ��=h��}����z&y�������u�h�k�Y[x��ڦ�K��G����j�� D��x#�;�����!��'��h�38a��88:���}O8�S������תW$ �P��z����x����6�Yd �� ��7�S�a��1�|o�_3H��cuʨ��e,�mX�	�:?j2U�d�u��A:.`�(Z��������H[IH�M?w��s����!��q~�����aU�\�9x��\���sn&��1PK�P��uW=�tn�y/L��o
�C��|����@Cѽ��&�,F��� �|�=0�8"r��2'��s:��nL��hi��9�Q�!˽��# &�a�'��,C��^��������VW-���~	G���犙+}��#�������#;s���i�Nf��E;�Jt�,�_�|���v�q�����b^��)Ķ'���-�l��/���@^�Bn��PahỨ�t�G&���Dp��`��_�׉B�Íh;7�E��������-ԩ�;z ��M��V"�N#cGmT@��r5a���|�)Mg�X��ǉ�G@�ɔ�X����t�t.a+��#�B�����l�4�["����L'|�d��x�)�i�?�{mLE�6n�hm��#��6�y���~Ȅ�oRo�&ߺB�����i���5#���+(����
�o��IHQ��5�Fb��q(8XwJ�(͊�&ʑ�c����얝���N�>Q �%m�'3��Q��D��a-��k�Jm������)��'��L!q��p~����ء��=4frrA��M�G߬E�� ~�F*�j�(R'�.ԑ̓�A*T��^w�����T���M	,d��`iP�K]�;�Ki��@P��)��рfJ����)
5i ��J��.9 y���l�����t��� ����[v&���k��)N���ExP�u��jh�Ԏ�q���Hr�� mʉ��;�ȸ�6�z�,iO�T*
�V�(�Ƕ�����!׽Q��{E��� ߷�W�3��$Eb��� �N�� a2t��-�BO����q��\	K#�<�����#���Is��7QA���r%늡��/׶M��b��ޖ��:N"�-+
��S�v��d�%��o��'���1�|$d<8�C�%�R:%Ę���^b�*���/��'���K�Io�@0e.�4jX��
(f��\f��6D���[��\U�m�x;�A��2J�B�C���jѾ(k���b��9$�����i	�-b��$)���QΏfآ�L�XN�E"����Dϛ��ǽ����\ַږF\i�ąs������O6@���3}�� �	����IxZe_ʸ�L�>�!H�x���^21�\f�|�R����������e� ǽ8��h���\:��%�{���O���e�}���8��5�w��Å]xĘ fJ��X⓻��*�S�:���]������6_����H�z+�k49��Q�M��ve���x��%��3�Wx�˿P1�xnr[�.����cf�J<�g��c�y���+W
,���$�)�>㺟�C�D���7�]E�����B4�&�� G����|����}
z����5� ]�},��y�E$�c�H6�5h����}B!���׾�F"+\��-���!W}�*��{�%ٵ�,/�+�x����m�8��Z���PЦ]����X�	�%b���?���0f�W��t(R$���r�:,���u�k�Y���q�ss)\�/��6	}_����RT.�GJ�}�޻���"�"���s�H�9��=����<��r��t\���P.�*ȩu�A��:��6�V[��.�>Cdy��&�+��y�lpN�U]���6YՆ�S8/�+Я�a�S��0�_D�re��K L�=�0[-x��F��A��q�v:�y���k3nh���q�8����W�ϗp����ᄫ�`�����c� ��}�&H��J���p�h��Nq��+�V�����K�06_�������WHc�GO��� =-^�Oc�l�)�fe�g<V��PcS���������p�Z2H+䵌dt�y4wͦ�F��c&)�Q�KT_K:�x\02�[O����S��w�h+�iB�Ug����;��� �t�#o���/����:���K���65J
�g9�V*��Lh�&���l�1��]0�H��c1U��+�[��K�WNȹs�,+Ԏ����O�c��y�~Q�ޫL�{����=)^c����)���\�:���Nl�8�����&�<�
�(T�xu��Gll&Gsw�.���{5�u�Iv�X#~厁���:N���4Q��ϐ|1U����Y����|Z֙�a>�2�v��Y�W�"8��L#�$�)NL�YM��l�_RD?���9���!G�V�P�%",q2Y���o�J	��sm����wmsr�_�(�Pf�1�l�1/�n��b�O(��'\Dtr��0�\�7�ݱ�EFx��*_��y$*5/�s��O���՗�u�Pz 1�[,~�T���3;s�<=3=��Kc��U�Q�9UhN�Bߐ�N!��}7'Yp1[���q3�Ri���I���8�6PaQ��k̞��ԑ3�H�A'^([N��ۀ/J�}�Eـ��ſ!�M^�z���U9(�����
V�]+W7�Fb��a%#�t�X|���ؒ���u��6zLӆ�d��ic-#R�g8��#��T�Lne���S��LV;A�M�i	�����,PU�O��a�#1o:*�<gB��Z��,�ǎ��Kœ�U�Q'�lN���y{1�_H��-w&�A�����f��3�Gn�WZ($�
34�7s���w".�+���\<؅g,p�ZꈧU��_0!�[=a�c������� 
��q?��v��MB� &y3G�r�L�����dX�t@q���go��%����.�v�\a�����%����W%�����C��&w�1г� ���k'�nld��{��Gs���}�X"gJ����of@��вt,z�'���2�|��1�Ճ�1���[�A^LڃgWS+ � �q�PfC�ߕ#+�է55T����jVG��5�=��O�	��$���r2���QJ:�N�~�+%������DZ���wӤM��W#Q�Bd].�D _~��M���� � AT�3�b涯�u��ᣎ�_��M�z9>��rhL�+$X)�, Y����p�jV�͇5�p��ͽ���̲�5�24�*�?����
����p]����$y{���f��e�SZYu���L�]���Z�6�h��]Y�6�b s%'W���w�d�-�]x$Xؒ�P���F;M�'���&Ð5,<_8z��|�U�؜}���z��fSP�/C�FvA���{�G��i���%ww��u>��h�ο:}�>7 �M�'v���e�׮� V`��N�S6����F0�"#S�\W%��G��R�|d�W�\K=[�_������L��˗L*���w�Q��:�N�C0�y��q���q=?�0.E�|�簮o"id�\�<�|��@�3U:&׫�r�,M~9���������Y�0+X�7�>�)C�{��IA+�շ^Y$-��Fn7ˈ��Gj}	纜%.���垊��(���x�cf0�����v�t�;d�Y&���ܣr���R=Y��fU �ƥ5ܥ��jx�Ww�:����`p�s��N�h#���߇#�,b=@��d����]�J��7��%������:��0�^�#��\DGI9�r��Hdy ؋=���^��"�4�cs��q���,�k�#��R����?���D����i?�"`z/��e�Ȳ�O�Fv��j0�i�+��k\�����ն��e�����c�*_T��uaɸ{9,�@�'�d!���h7�i���M�����q�Rb$s6�eX�fiw+w����rgdBF��D��"����u���h���(mm
sX֖�ws���@m�1s���eC��j�fԩ�7夸�!^D����!7��1���E#�BOLtS�#�D�h�d��ɒ� K�f��%a@Ȏ����G���B�W^��X��`}@�ׯk˝����"9��DP1�{E�	8;��~HY��`�'���(�0'�IW9R��/��&��e+�H<����[j�!좫��T��s��B�Q ~H俜����u�k�PN�E�@]x��#G���}=��9(wO/S�ߵϯHUlN~?g�3ר����s,�x#a��|�v��|�l�������;��� ��,�ѧ��=��Ӗk�Ż�U������X���&(�02to�q:� d��R�/7:�:��LD�QB>]�@,�����K�ATڶ�����!�T7��#ё�C2���,,�4�����Oik΄�jj���U^'��y��x�7�2�Gv$��sr����P?_���z���;i }	��j�K4k�[|�J�/À@o���G�#�W��Bqu�d�?������S���n`!I^A���쑥!�k(����z$�I��� _�>�����?���7���!�Ǵ 7������4�fpxO��_��㒥||��_ǡ�7^S�s1��L�h�)��άB�S?��4,Z:���._b>a�=���[D����:�l��{a��(T�l���~rƤ��r�sZS�����4ի�U� ���Dqs�XzSkB9mĽ�����r�s�����M��=
��u�Q4�;f(e@�.��\ ��JPÎ2B��P�"˵��h�3;�������t)[�n��E�:��K4"&&Ӓ���_]$GD�n��3P���{"]�B�͍����	 H&����>��S�B�#xڥ�暴�7s��B��](H��9g��՛o����Cߤ��qo��K�K�:b�=C1�+�P@P�!
�`�>��Y� �N�'a��SL��/|�Ā�&^�o��"i��i�ò����<���V���6��� �?����g�Sv�wħ���H>t�.$��� �2̒l��J����%���v~�������"{�f'�E�oR��G��x?N�]<v5��"R�6��(x;�)��v����3U����0_=��贴d�2mrr��tx��o�P��!��|�[�J��!Ux~����Ӟ�W���R)w���qG~�� [��wX윤~;���+��iHK�5��,���'1ܧ\��/�ԫt1�7�e1�]�BJh�t/ �*t��9��::��7�>]2ze�nH��Es��n��,=޵#DE��Բ����3�D�ش�M�7���sZ�҇4� �Cp���4��[�$�g��є5ȸ������"tR��M���5�C����66Ĝ�s��I�����e�ZT�	sI!6��5�MH�G�A?�47 R٧�'p��$��T䚣Pߏ�u�a�av
ȥ�aS�"�ooj�y:g]П�{�<��OVIW������,3�_�>0tuRp ��z8��-w��>�W� \]��x\J��n�m>�m~g��k�x=)�����\��F�*W5�>��;��kiӽ�M#ю�O��r��B1v���.G�-2��8��ϵ����V{����_6��#�K���(�uX��≢��R��6�۵8� �o��c���ع��T�e��B6���C����l�Z����>���p.h�na��n�#I �wc[�+��ַΗ�#"�TM0u�pX��n����3X�M}�%���_ml3ܷ��jt<Y�8%����M�������%��}&|�6��3E��ȸU@�8�~�� )d�W�i���@T�RRJ1qD�Z�D���Agݫ%ـ��N��Q=+��ey��+|!��N�r�Gq��LD�-�u��`�ﺃ�W}l&/m|�kǠ'�Ms봱���ߌ�'�.�9�N���TE��\@�s(�A����uRC�F�,X�'���x�x�=�]������`� �J�^�+S�����ќ�� �kE�����#��R�|XN�������DYɩ��R���s��qK���E��$6n5�+�tuė�o�	�0A�T��#k�c
!���h巟�9k(O��<?d7Y��ZA2=�ҾL�TrN)�.	d=o�#�0��g���t,��k͟�M����]���Xo�/�� ���*��Eu�m�L+,D��YHG�+��_T\���=��Axu�� U�e�ףP�O��W��3��>NE����V���v��ws�z�!�䛋d�KJ���Ū��))�[�>�;�#�����0�ݵ����G���7�f�&A�q�e�x�Ê5J��d�M�R�h��h<�^�`�9
$X�9WqJA��
o�[�:\�>��=���w��j^]�`�E�s`���i����>�@ �G��r�tRz�ǁ��q7*X<�|/Y^˄'�w��?*t����-	����\����7��+�)S�v�D�I}&�}u�
�u\���Ι����YF�Å�j��_��wmv���Ӆ���7�nsG*�ÿJ#�]5� ����̋������y��܋������ZmS
��(���DMD���Z�q��� ��D�v�qG�AK� Dv5K�(�:W�4�Ğ9(<����J�`~zT<f�٪̞ڳ�I��t� ���z�0o���O�Z�ݐ� )Y���|,�z}����}A��9"�\.%l��a��.;�B��;��0m�_�n��4W�V���(�����oRh)P1�-��w'1�˲��$�����f��]�I�Q� ���p,y���!y�ɵ�©B��TG]DV�UDp{#'�l��z^`7�����JVC��r�K�NE�>[]���٨�OB�'){��7�B�����u�_;�͵�x8TہY� L��H����!. 6h��C���7���P�»����V����&��׽{v��������<��JQ8�R"Q��\3F����@^��x�"�nh[�W�<��J��nO^af>��!��ɫo�h��h8���6���6���
Xz���h�)����'�@��F��ã�x���܄�>�����@�ȵ)`�-�[вtd�$x�(n���JU��pr@���|��p�O+�:�����50�P��p�=U������Vgǰ�7Z�i�!`t>=�l`c�_������$5Y��Z|�������QPs��v~J���dl}������qg�ў��������\����r��D<��~寁E"�����zL3 �+Y�Q��^PZ#�4��X3ܜ��~�i��z	��Ĕ�}+����DEpW!�e�����sXeu=�L�pR[ e�L�w�	�LT���rU�Õ����un(6	�:2��u���bq�W�tM�O	��`G��V�FI����X����ia ׈�\�FiCd[����J���>���P�L/�@��Tt�{j��7_P�{���?_p �[&��AL�	���D��G:׻�r��{cΠ�HCJ����p��X
_J4L�8�3^C	������¼$�������zLq"
e�m�����#R^R�y��Z�z�/g�F��ȇ���Gtl���u�ê��g��V/�%�.vw}�V��[�9�US��P7�MT�{T???�ϟ'�K�M֩����������><��Ψx/UKK����Y ��ٖ�ej�&�C���Z,L�T�J�5�jeDx�5u����=uPo�Gz�E��fR���8�U��?Y�E�c��-͖�-t`����cx�'i��:��@�+��Ş
P�bl��g�`�wo�TZ���Ey��	�e�3G�֡�����z�P���n�f+>��Ľʺ�{ҊuRb��R���${t��2��%�Սf��!�/�������N&����j�Ѩu��RHʭ>v5����*�h�M4�64Lo����޲$v��}5UU�_�n��h���.������2������]�~�E���U�T���2(T�j�3����R�$&�����'��*'|�j���)XcSw�S7��sEi!&�"��fD»��3�?��G�>��$�s�����֮~����%
+yu��'e���/��1gA�pl�w��AΈt�C�\�) b�c���%a�$�Ps���+n?�/y5j�v�,\�B�L5W*����@i�g�����Y	^;&���7�4>F/���L��م#�@�������g� C�ND�ujRA�ܣ~�h��]���4�}Hq���rI~B�^�?�R�--9l����-�X� L�'W��ii���u�Y�U���첵�ާhk?m��h�?� ��(��q���/	��b�����͌,�Q(ԡ�M��T�kᡟ��r~�T�f�������'t��C��6J�g�Ot� �`s���Qrh.�R)��ÓRq���* [��p�}^V���R�L}��I������E1�~�m�Fׯ}���0���p����Hg�*�UW)�{ �Q�_�E		�Ѩ�E���+����-\���Lk#�G�c�..2}��ƌOʶ�N���,��]��J��=����0Ҍ�6������E��򋌻���>��a [qI����	�J!u	�c�
jk_[XXܳt�pw?2/#�v��n�fxLqSSx���`��� �НM��#k�V��-aH��Gw���<�ua��p�>�����Mr�)��s�mJ�}�:����+y����x��l� �E���Z������
��Þ������K���KA
��Υ������9���?��(�L��T��W�zS�L�c�+���ݡah-Ǽ������҄��p���?����S��1�ݦTFDD0��8x�����䣋�*�L-MMI���ݶ'3�� ���BL�~hJ�Ib������/ظԻ�v�ad%=l�hy�.������U3��7{M�(!�/3��	����#!�IHH)�K|��=��_��#�?5)�ݯ�y�1ݘ�?.�^�&����[3[�h�_���T��?X���4ǃSʈr��5������k�	d��m���~�t��"1��}"��V�*�4�f�ph�ۗ��¦&B�H�F�gn�J�ާ���$��eR��9/����^>���N=��,W�)e��\��O3`�7^���Q�gs���71<+�3K�jnNJHH�ʔ6&��yUTB&��
[w�P�K�[ܙn��lK�����ޚ���M8��6���S��^U�.�ض��+�\���3Nh���<�s����ò*x7�
��ni+�ld=���t��. fҼ����F���z1�fc��<�����|̯=��"{�t�@AK���ʑ�q:؄<�k�#���:�1�gG���vn/hG���|�v����7o�j� �b3l4T�qmlj���)��Q1�IC'|�{T��l �Vr��|��O��ù��_�dCX�=���h}�=5���/{4�7�9�2)�U�I�^����m� 6��}6������j��z�j�ܛ��)�G���l��+%n����ݖB=إz�(ү�*{��_<�@UÙ|���ꐉH��p�~��a���YϹ��j $��,�6�_��Z��۸��du��;�C*6s�
23�V��TA{�J}P�*o�Ǟ�2:�"�Ɖ��LG�&#�Q��A�K���q�m��_���r��$����UGUjk]Uz��T$i �.��=b�MHPFGP�j��zQ}�������>@���9~KKz+Y��l4���W0�ˮO�fkf�1�w�!�%�k�?��,����T{�����>�F�|"�I�Ǚ��T��=����:jP4�4!���׃3[���ԺMa�����Ɨ���b_��`��;��]P8t�W�d�.���g��oE�� �_p�y�5]F���+��2�Au�
�h2�����ǘ�A�AJi�
�'��Ds�tv�.��47�\�����a3�� ;ۛ ����~r�3�H��jk���a�hن�*��@R�:�6J��7Z��?��B�����,�;O���R9ѵyQ�9��g��|^	q�x����m�nN����#��3xd��>|Ԟ�����9�0�2C�u�RͅR����<F�;>$����8|9n��.o1��ė+�b{>��]õ�QLX_��_�D�!%ل�2�՞�IH8w%��['``6�i�r�Os�o÷= �0��ځ+W��u/v�4��<���<q��9�L2�@Ӣ^Y�	M�ظ�z�&SK8��J��/�@�	���c��J9���ˤ�3�h��c��^0^o��t�Lax�o�t�W��S��y����ښᾼ���H�7�T�{�CBA
����A���m������8�(�aZ9�*��H2����ۄ�t4�I��1��9�y�X��2o�����[��M[l�u聏[ZZ�KKK33�[A�	|Hf5�fhꈫ�����*�!�Io��G���ׯ��0��)�?'^cb4W�8棦���
%�s9\rU��P�LǢ��
�xsJ;"d3�5[��kFF���j������ls��B΂4�}ZEDx�����ʧ\V�3��>����R�{�%� �^e���0�F �0���0@���i1�8yD	~��G��9���ō���77?����8�kQPs8����ʢLw�����:?:���4����׵DFS-<<�Q[�����nB.q"W��o>����=�N�{����O�Ne1�a�`�>a�e��7e�2�f^�k�[�&v+�ǳ���zhO�������SRV���]][B��/џ��t��񵴂�@--�k^��NC9��%���=��^ߨ���x�u=HHT^�b� 61�m(3ȧ'�33K��4�Gh�
`��ɖA������w���\��>�I�.WK�ҽ�G.yJ.�t�qa��:��Z�����V�7WWs��O��ꅍ4����"O��!���-�뱖Fx��{��C�����,@�y�J_�&U���3]a����VX��Y'���i;�nL&gd��Z�aQ�[�'O&���,�;H�g<��'�� �c1��7�=�	�������-�H������xS�m����B̓�1��+�tS�)����MMj�rB��^ý
�}rX�'����7�L���̟��~�dX�<U����4�:Uw_ʙ4����{��t�΅���_4A,u`�"��h������T����"���jt� 蒦��x��cjo"�C�Xd���`�	I�ć���OOÑ��/\4��a�B��J�j%����c4� �"ZA�ܾ��L���`E�h���+�?������޳�����7�������Ip�6lQ֛�����>7�u:�i��z�Q�"�/E�|+̇m���"Z�����D��j\��[�3�ڎ� ������{�_L�� YP�j�FӲ4l�$($	l�vqE�DX�A�:�i:doo��rm<Z�∆q���ǂϲKV
�TUe�6V�&4_K?Z����=`#w�ɛ�6M)�^,�rv;�{��@����� �w>������\������ �
	���'ΐ�w�O�L~\ C�%f��®���j�lT�Ք���dz�	7��,ͅ|vf2���e�;<��{c�5,<���Ϩ�NH��"�<��3�}���D��q@�fm����xgV��˸�Jb<#Z�RR�Gl�D��{W�f
	�^H�I��?�=�A�~����Z�r�;�]�)o�la+Z����ߢ���4�w�\��AA�q�c~AACX#GR��|vFA�oSv1x)�Q�V���J|>���>zm�p�op�C4ȓ�@:V��f�k��垹�����]�G ��3k2[����n3Z��~	�Y7w�k��t�u��X
>���ޚ����Y�8%���zݷ{�x,���= � ��D�\jx �\�ء.�M����;�R�'���^<q	,�V~�0�a����M���Q�d�܁ˮ��`0�yJ8 j`.  Xee�-tu�G�,��;1�
KƱ�`�i���.p؞�-��k���N�e�0on��N��:; �=
z��rv�{�Ϋ��)��h ,#�J�?�r?�]H���1�jQQ�����C`S�����ͳ��N�h@M�r�pwxԡ54�m]P�����F	�I���w�､���<�/�q�ŏx �S��1����z�H˷����>�T4^�x��/�m���H����֔@�u)��6�#�2Y������������t��ƭ�M�R7$dTv�R:$��I��{(!�ށ���k7|j�W����/�qUQR����2)M�����'�8���b3X�=Z~����:�FVV�#�<�G���M&>�{��|���>�:��u�������i�O�&m�|�Ӯ� ���{�!��VJ/ҩ`�]R�@���+����उw�5�� ~��Gj�кm,@pH��u�KK��l�2ž?�ʅ�B���~BB��H�W�!$���� h9U>�h:*����֭[3ǳMo��r�����u������ ݴ���m/=&���H�,�n�a���!�+;a���-9�HRAoVߎg+8	�- ���[��x �PZ��B$�A}���%dB)�.h>!x��Ѱ���>�����<>o�s���<R[�����f?���Xo�h�r(������K�J񫏥N���T`�C��4�hdO0�ؙ����6�{��t@TopNX"�&:�}�5si��t\	��%�c�UX�:ލXJ���F�~�=����\3܁��4�e8���jdk7^�AF�����ϳe=}�t	��@��Դ���<\+*	���ǹe�v=�NI�=�?��|N��d3���m8!��@^zS8ݿ��*����V\@�i-���0  �#�!�Z7�ӵ��҃V{<��Ȅ_��HUU����Wh�?��t� [��jLw�׳�s`bem[/�9N��;-y��m��E	��
�������[]��W�d	D,H�KMJ�Z��T��1:ȦN����@���C�Wa��z= 9nS�������
"�H�,�h��t�E���h�p`ݿ��v��=�6��P�e�+�Y�Ӎ�_y�\`��
]��WCdx����st��DE,���*B��X@IP�Ca����@6@o+��ӏ��*='g�p��@	655Y
Ս�s*�/Tު �`�a%��tX_v	�������e�W�|5\�<z�<J����H�oc� � 0�.G�8��p����z�G��/1(�z?��?��ش;t�k�X6N����m���$��;�^'I���Rᵶղ�CO� ���0��G���A�{���� O����V2��W3�[C�\�Nk�?��DaS��>��E�s��-`��(AZfz�t1�oj��c8�3V��z���'_Ց�<����B�}w\��7���"�Y3�������W˅?�$�Ē�'�C|�8/�@��t�o\ٴ�#� �7@B�#��ҒOw��+%1{���\û0�����.A-ű=�Yr|U���GzL�d'y�%�o�F������Q`��.�B1�+h�e)f,��}Ŋ�fKj]n�w���V��$B��7�k�o3 ���"8�?�& BN�h	�� �X�@������=A�Sʮ7��+N5�gi��9K�X�W��{0��U�.w�O�����y�o.�~���f�2�h�9����pߋ�����B9��\a����;�v���<�д�	�!g�~E]���꽃U�z�TX�:#%e5�O���S�U�	��?��a�|k�l����4�����w�x�w���j����C��V.�X�k8�ి�������ғ�"�䫃^g�o}�/:��7D���Z��vK�G��&�g��� ^Uu � 	!Bؒ���p�"���K�vY� �:=��_w^�xj���Uś��9g��{}��J�k�n�QH�bE�Q p8iF�X����p�c��|1�<�����s�Z���ƥi)�	j-6�x<�� U�wsSt��mM� !�ޭ���2 �7�?�⊏�u��_��։l��*Ӝ%� ��N��w��?֚��������2�QQ�For}�|�T�� p�W߫ �)d�ƕ}8�*̛���4g�����V���+M��sZ|��_j�G3?
�y�=����'4���l������(Nʟ�o��qڢS6'�����η^�u*)w\�ⶻ��k {��+�}<R;��Ԇ0�m]=as�Ƥ��/�'�v�r����[�R�S()�z;����g T���ٳƼp]��g��2Iʋ�b�A��+���~�j��A,�ȪW�dXL/�$�F9*粊����d���Q~���Y��E�����IitluS�c4�:x�6l\�=��iQg���ɛ���ϱjNLG�4��a3}Τ�H�Y���\���۫||����{�Fi�؍�ʹi���N��7���z��Dn���	���Q1�DJHCj�R}��w$+�E�U�}���m�:"趶^=$드w��˪�
!�M$���3��1���Uc#�Bw$,R�uyS���C����:������	�^�KTrk:6W��:_,_c�-*����ob�+��nt�)�.!yG�s�}�4��*}���lI��#��S;�M�I��#h:���]L|c �����))�U5���ϡ鎊�ec��*	��R+�n]�+73_��Xr�0�[��x���H���T���S1�#)I�G����H�x�1^������-�)��߿_VWP+���\fw�X���"����*�eT����J������?�^w�a%t�ˑ߆-��TF{�2�i��J~;f�n���J��QT�yR�|͞G���q�\V����l�����*?j�|�P&�]����1�ʑ������d�B�ŉUHc�D�]�n��<���
V�w�hVXIu��'`���rA�N�d�A܎���Φ��j蔥�dՉ�C>���=ΚwX���bb"��%���>�lm,f�`<��k61Y���
 �b�"�J�Od��LM9/��/۱E���֫�'�D6��{���Ɣ�둧�iw-����o^.HB�����O���	<�T)D%,oV����Ϗ*̛vU�q�IB�pYh	Ra�s�j�E���D��US�J�����CW5�U��`�*Jj(:(c��-��=n��<I��a=�Hb":��\oG-|űvƅ���"���x�I��J������) #����@ʬ�]���W Im�@d��GK�I �>/���\ʮz���潵m�i�{mU�Xy��$kE�~�'2A2�&I�v$ջ�.'�Ur�!^��Tgǧ�pJ1ܿ�JC��q�+�OTd �	�I��zM���(s���^�;�3�~7�1m�]�/ 8 ��`�($ݚ�e�(v��5����e¬	��Ud��W��>�*���Ԃm>�:�$��Dӓ6fV�y�s8�N��s�Xg����-���UMVH`�9��5�A@�_6��WF���t�r�-Y�oV���V.	��>FxA�*Ӯ��T�I�'�n��A%T:��}�J"���i�6�d���3�[)�����D�a�e��f��}�rkn��%�L�����S�\WہM���R1��H��?*ts�ޭ���`���#Q����|�Iu���Qy|՝�]O�{������E���&@Ⱥ��X�	]�%�9<��x  ����%�H�dZ�.�,�|���e��������z���9`A��v���Tb>;�%�M��a�o$`c
��1U1� ���aS��d��0�<�� ���Pt��މ!�I��q�&�s۰TN���pk�mƻ��3h,�s;|�ӱԠ&׊����T�Jy�Y���_�j��8��U�Z_�.;ݱ��t��B �yRڴ�Zρ%n����Cʶ���0��17-��H^L�tʾ
�-~w,�2���(�ex��3J{E�_p�:�����$���� f8��!p���N�W[`�^B��C%�i�~���M�J�4J�F狩��6�Њ�C���	��BY�kg����<%�
���"�M:��HAp�ՌP��{��â����&�#�wY�"*�3K�V�����^[|m��<�z��%�8b.����ԢDx�/��y���,2+�p�����
d����Ti�46/ ��v��{��]���I���5i9Ǭ �u�����h2	�Q��V��p������1��JQa�+*Y9�(n�jn}s�-ہ�հ���.{��Y�²�MBbD�a�V��9 %N஭�/��1�*�mv>������m�\����O�{gݐq@���嘃xvҞ�V��9��/'�s <��$�� �,�1���`��T1������=/(;�Rr��@� 5��g2?� ���'V��(�ۼwI�x�(#�A�:0ȹ=X�kjA�v��@ �`���������y���(������k�.�UV��$_�������o ����Z�e!�pXv^t��_�Rl�}�^�>���CTxT$�ы/����loC� ����y��w�rvռme��TTp�&J1���"�U��*=�j��|�V�C���~}����,��pl3�+�'��A�݁-Z�sxW��R���n`&��[�o-��b���::���_��v���B ͽ��RM��D�e"�\�Gd��r�_��R�*Q�/�Ի)��v����D�ń@��g8�iL'�����3ޗC6�1*"!�3ޭK�8*Ո�'�=��u�"����ZA%a�m*z�������m��W�F��R73��X�N��|$Ǟ�o6�'�4�������daV�x�6L?�,�vv#�A��u���d-O��`���lR�!u��x�?���mЦF�`k��U���(����m���.&5��
�ӻ� ����6�|��		���~ܮ`t|�7�]�ݜ�f!7
���Md� (� ��(סuh��dw�0��$�|��N9q��m�������)P��|�]U����[��B�9���c�F�x'��y/���4���L qm�cl���r���� �:�B�=�E��u5�y�lכ�g��5uH��䌍Ns�p��w���Xp�M�����DԉR�O_�<EeF��t?�]�q C�����ܐ�T��T��S��B`�~#y��փGvIv2q���Ͻ1�9#�������l� ��>b�B�b?�4q(��ѣ���bf9g �+�����\aU|1-�U*��f>~�m<�I?�G�3�]�4/�=p�j�ƨ+ �ms���?�y��t �<T3�?&�r��N�����B��t�������L�'��x�2�����T
*�gY=uӓ�w��t�-=��c| �0����us~t���vX��
��.��]{X�h��	K���m����5P�w��e�"�yᑔ@��p��̌{;�?�:��9��I��Oa��O�t�,@gN�y�=�')����:2W�xAu�	��b  �R]�|�4V9m���0��iU9 n5
06Wt�5�����}㔖T�	^����+@_;�A��B�`]iG%� �EA2a�03Hs_[���EE����C�ԂkfW�`�q8B��S({9cG߸�v��2���TYS{5��y��!���[Z�����*�Yx��+�~U�H)1���}G4����ҹNiW��V���Y�?O?��� ꀦWs !?�ce�ܭ�z*��m�t_�_�P���/"-:�Ż̎����R�RVl���I�a�]�����W `9�
��Z c(�l:ꪊ|�*�D�P��H������D�;�b�+�:6�h�� !Vt����OO.��4J>����{lx�@H������mۧ�O�p��M1���&ٔ��5��G�a��G�d��
1��os��l\�_ف�#��\k�P����5�~����|�y�jN��+�G�ē��V�X�$*.,��	(n��Y�V\ͳ��V���
�1�/�����q88���%��%�	���Q�e������	"��`�ײ2]dwmӵػS-��J�B�*cˡ܀�d���Tk��
�@QxCϑ��L��~�ygIM�T�K8�3JCq�Р�M�i($_j�JjI[73�~���TJ�"��C+Edv޳aq �DyҌ��jf�!��=���-f�cD�tN�����j��yy���#������<�����d�v���|Q��%�"����S���{슋�D�{!%w^�Hu1�����I
k�n�T�.]B�u��,�`M()kˣK�IE��e�lޱ5�V��.�຺"�c[v�
��@,�����>?JT?bk3��BPC#ԵVn�0Z��#����H������6��w��Z������~@4I��b.�H�A�,Ѡ����;�����k�(��m����,��{l����^�DE�dEQ�� �D{�,���pBX�h�nbG�iy���x���+�]�c"�M���E����_�Xp����#�l���KEd �I���f}��>9�@�m;����}kT/��H������66�LdIjʽ��:
ʈn��n�fT�ӌX���Z˹�)���GʗB������jwkӵ�%�r�9�r�J��Ñ;��5�v�,BH�F�����P��cr51�䘤1!3�q���9J�J�������z=����|���E�a�ϲ93���o���7�<�(Z*&GI��	Z�"��Ⲷ��Ɖ!$����Ln�ir�K(���g5f�u�:��dx �-�o�a��3.�X�g�V����A�Lzv"q���k�F���͚�������틏�V�!�J���� ��3���p��m��(ź|��
 �y�PYN%!������T�*� �AzsV\�:
����.��uS�=��� ����X&#f=v��?��]7\���-�� �;$q�5O�Ӱ�7��u�=ֻ�oj���D�ֻ����U���q5]���eF���ЪB��a��o���2�
��e����`R��
�0��Ԙ��m���Wz(gh=52ڌ��3�ܢ�����jf���E�P�Q`~<�m���9������O1!��;d�ؿq[F�IQ��;x�bm��&J+���<��w���q8qw�X�o_á%
#`
O���R'�Dt̥/	-�{��{��wͺ ��55�4}���U��Z�DJ����\�S���,�PU��d�w�.��;�E�W�)�s����!���xW���&�C-� ag�B
��uuu�Q,�AZŪ�_M:`�!�b(}�i����_����-�)%�����"Nm^C��B��(3mg�EH�։�ȕ�]�}cH�D��7G:l�ɶjO� ��C���8|����]�e<���jPTP1�ȯ�U�k��t��c#��	aM�z�e��'I`v#CI`Z3v�ͬ/
���+�y	��\��)�Yj�{�Kg��<��.�����eߋ�>��������.�Y�Q_H�k`�'(�s4d�$c�c�y�*Q��8�U�y�F��H�h ��g�D���i�/�Z�`BƖ�����^~ ���-3oBid���\������������%�b"}Ws�:��,S�e8�if*�کur�㤉=j5��}�� -X9�- �:wp���=�=��� �c�fB�P��k�f]l���H|t�lHI�5�&1 �덂�p6�Zv��W��;^;��ߞ��2���<���v��.�R�+q~�A���2��(�Shv��W+��	3�ɰx�7�E��������o�����:���wW8�Y����>�{\�7���`BE���hN z��/�
��A�ř������~͌������+���T��+��L9�<ջ|h��.)w�@�Ov��H�k``|��w��L/�w;��/je�P�˛�*nʮ�����!N�S0�5͐GV���z�e�R���?ΨU�q��0B�JD'��Re�xD�]�y'�||��*��`U�w���jT�U���w|4.q�̢�8�3�����u����K��z�o��T��c��B�l�/��,�0��r"���.j3|֏��,;E��Ht	�ZL�+�W�34�o�?��M��>j�8���&�~��Wz��VM�y�T��yE��;�v�"{��c�
q�a��=^Z�)�f���0X�Ҝ|�wIΠ�!���-����<B$�(Q��kD�E��;L�<c-U|RQ�k��~�]���y�}8G]���5C�U3��� `{2�[b�����@�{d��"��5@&Xc����Ŷ���EW��Äԟ@�`�$��Jm�[c���RNn���#]nfXؙ��7�ݍ�Ȅ�P}����aREW6B=�:"�A}ogb��&^>G�_�g1���C�����b���.�`4:0��w���K�dA�0�l�q�*�	a%H������X��͙�~��\.�{��69��1�J'd�w��.�B�T���z�?Ӫ��d��Rj�[����x��eL�D�(�!ۯ�R8u����@MM�M��g�C*1}h b�W�k�n=I]3Ò�0�;��ܔh��s#��Z\j��`���F�dQ�S؂����2�U"g�X��w �f��P��<몦���� .�!���W��=]���mQ�;I�if��=�r	�t��S��%��5W�pf�p�|Mb"IEE����Ţ"e
YVDȘ��w���h]j�qh�=F�ᕌI���`�|�v@�������;�|��oB�vkR� *�p)��{.j�^B��_��u����/6;�����l�ҍ�
*�Z�u��p��EX��!3,�������͙>I\j	*T������b%�r�݊��N<�龓X����G F�^�/XW���3?�%��3���o&�k�c+��-�(/2�3;�E��{�f����l���{?yt���Ec`���8�	l\Z�8Ԯp"����zz
'��V!���IaS?<�7�sQ���ٔ��4��6J�5o��O���Q�Te�&pB�����(?P"�;E���A�U$7
�r��1cB�J�|��ZJ��ƨ�g�U[�]��D���GC]��}˂53I�j�h����S���}��ե�_Q,˽5���4�vƚ˂A� Ȼ���hRY"�1h�z<�=PӀC������g�$1WhY�`oNF�D�e籣���W�`7�]_$:`!�Ҧ~tm{�Ȅ���?or���$5�9f}�Ԍ�j�6����&A|����p�cհł�S�*soR�8���$�>!5d,���қ�������������z�\�Բ5<o��s��WU��F�X���-c|�8�&�L���cz��D�}l�|���u�mRLG�]��"��8��ΜW�����H�ƭ�K�$9�q��x�.����


�`wU+A�c@��I��������+���;�koJ�<-�TO$.�4�W��@�ov��P$s�;k�d0'N\,�\���#oH.�*n�3�X���PB<f�yk���j���R�9�A�� |�h�Z6-�v4��`��i�Ԡ�}(�;�I@k��� ��+*Ğc�vy�?n��格 ����)Я0�%���x�9^���ΰt��ݝcMփ�H}�_���P�ߡ~%��q�r�{>��ק��&E�����M�gI��o[j i���3�p���������Y��l���W����j#�w�����"zچ�|7�2�Y��p���=Nm�TNkl��J�O59q���>"i�6�Ȼ�����_H���Y��)x�づ1EEEOR�DEt��"�#

d���c>1�[y� �4֠����x��m�Jζ��tݞ�����A�(
���垯��ԡ���'�o#	�"D�O�X�ց�@�3�^^a�Ι,A�����z��AF6��̠�2����������D�F_��B��Z�'9���>+�"^1��K�Y',������V�}��Y��P`c^ί�V��U�nJm��sR`＄Z-mE}$��W(�cղ��R��F����HO�P����W'%�P�(��6�.��' ����j��H�͎���>i������L5�y�B��| $�̐����"W���u��'���"� Z»���͡��|:A|B68�J_Bt��F�z�+�Ȁ�5�����#&��_��G�Emp3�kí�%��(q��2�&��^�v{����#s��RKp�0S�x���I�x��Pe�_>h_Wx�1 ���\jբE��e���ٰ36u�<�{1-j����/RA�4��<��&a.�XQ�}�I/������idvN�z&�y{JA2��6�|�/e���VNK��˸���Uoq�tc�Y���w�{���B�lc�ߩ��;ķ��'ik+�?��T���e�.T~[D�ci��P�����B�w���.�L.X��f��VP�Y���ҁW�^�2O2:_�����b�d��_���5�����`��a�T�sB�z� #��vFh$���2PJ$�}�&�!���?.߱�-��3�0P�`>c�K�M��vJ���I܏��9���{�#�pY����	97�	�m�m)���
�61�nM}��Y�5����Ȭc:{��߯3:M�](��o����������c�$src�%a�]>����9�W�������̕�і[Y�J�(G��R�u�z�+U�)���
�T�k�tT�ؚk�U9�m?M��l����a��ߏ��M-�bt���ܕ ���P�B}{g�5k7ؔ��������Z���a��f��Y��δ��L���o�g����Z�P[C�{�OhvTK0�o����f��9c���/s���Hf&�%W�9;��@���e��2�[z��&Շ2v��_F�J���>���R�_fQ���>���7�jU�aB�8�W�ςw-j�]���緉D*Ͳ�c�q�	D�6�{5��WUq��i,9̈́�b�1�3m�)`>J�BG������_��*/�X�ۃy����_�/���= wQ�	`�QZ�zM�!h���X��C_"<��zt ������>�i��N��1u�b�/xB�@Ň3~z��� ��g�^��3I�Z����ޣv0���#l�(��	 ����J�$�'���Ы�Pb(�f"�lJ�o��y��(+�xI1�h�l�V�CEㆢ�:Nė�J�h�ʻʅ��V�����eW���W!2�W�g���]θ�򙵈�;��>��n���
�o����}��!1֐f_�͇@ߣFf�7���]�J��u}2Ȋ�#h5�<�1�Ȍ�*
y9���C�{{�3�f�X�|O���{�E���{�������B��H��q� 7޽#�L�&��Feff���?��+ ��F�R��/zx�r�ơ�MA=�v�@����a�M���ϊ�k&�^�ym�y0���p��N�0��d&�8���J�|��Q�%� �	U7nn<29A�|���(�$ �K$�XGC?{�� ��V9���類�j���F�K[�ں	r3O��fOԋT���ܒ��z���>��]��t�TN�CQ�{r�tR�kp�w�����p6� ����k~,��}��)��B�̛�h�jg����1��W[r����m3�n/?��֟���	�h��d�i{)��R��@�!~fo�;g8��Ԫ��D�����E��z	L�ލ�u��jX�`��6TK�5`S��8���Z�Zc[Fڨ$�0F�v����""�͟i�i&E�@|�OQ��T�Dqaᡁ6�fC�z�	V!�R@����$g`ou�])^Dg1�>:��B�aW��f_>'Q3��[��������Hx��f����GPd�����h���dO����bn�K@RQ�'��K6�u�Du���zǆA�̲�SW��EE�uG����W���w]b/�B��sD4����~�u�mL$�W����T����+���H�9�]�z;�'!0/`� d^����~=���
$�!�?��u����JX�%��U�M���E��'�T�.((Hq����eRAd��#��5�:�v.�O�35+�g�G�rZv_��?&��f�x_'VSST��슰�Ś��~���$���y��$�8�39�34Bb�}�����t�� ��Դ��r��P����W����]�3��O&\��G�mukTb�m�e���3�A#��p� )Y�a Yf���l�����.��J��KE���&0��&Ǒ8!��iU+?t5�N�����WuS���|v�۠P0u��Ӆ���w����0*�ӈ.��3^
r<�6���`��|df�& �!�|K:+���� ��*QA�w�b9˼.�W�1Rq5Z`L�1�Z ک�(�<����+�Oa�iY!��=
{ޥ���i������&;6ႏӲ�`S��
����A|��Ǐ[?C`cL"6����	����NG/��Ŝ�K�B�X4��[�b��xR�V�\���=3�������4�����6�_WS��B��=������? ���/TP�|H��	�����<Ƚc=)Z;!��#��/��	^	M����$��KK@s�	��=����t�2�y:Ř�)x�|�����`���w��p?(�m_���-��ei��E��Pݙ������0n��pM��p��&�hCb7�=��u�����#�1�?����]���C��2�e.�3�C �CW�t��>��T����q�;����)�֖�h�^i3���O��ai�LA�5؃4���Ǆ�,=9$=)�\�����fg��i�'@�x@K�zR���y�5ԗ��k�d�XP�?��5j�|G� SN^��5KkoQc�N� � Q��DI�&�0x���@�悠S���0"QTnn��,��R͡β��֘�/�)�����X՜� �o��@���Eҧ��	gmg�g]xy�]�}�u� �?�3�ʳP�\�xc���%��8AƳ�r<V�j%�W��I�'\J�{�`�o^,�y�Y%��c}F�Dn�nn��i ��u�Kq�fѕ�nh��Z,\��8�ۑ���CWɚZyOZ�ƴ�jp��>�����x#
���B�S<�NA���|���^����J�`T?����U)��2�IIT��p#���*��S0)�	{|aa��		뀑(c��Y�eP Uҥmm�pc� r�|��s:��K���J���|q�`*t�/wġ��[��R!�GЌ	����*��Z��o�R������������.��D���S�r��"D���x��z��Pܔã+������5Լ��J�����輓�?���%عI�[�wKy-z@O3[�	� ��'62̗�b:�(f������ܧH�p'�&ת��Ec���`�H%(h�NÝ&'���o��*%2?����B��l}�{�	Ϫ�>��W6�U��I|�h�ބ[T�f���쫅<j�����4�����B)���Ӳ���r�Cd��t�O��P��F�r�S��l�GC��< 0j���|f�k���c���}�%�f������1ؖAmU]����w���׺��x�ic�ȻQ>Y��}�E
t�ahy�X'�˭��8��Ԫ��-��B� �ڋ��v��?f^�{�u��=����پ�xj=���ly�`�C���;����v��	g�~������55��/���71f8�Y�mP W���E�ʮ���N�޶���X����*5�%�ͳõ ��F��0�m'"��A��������ҪT �w?�t��Z�>��[/��<Q_�S�[��_��U��)U�3:7,�X��7�bNY}�}�?��g�i�u���jps�g��%-�!�����d�t�dP����_����Q�vf^���%����W�*��M9�e��pvy�X!�|H�ڱ�m\(�1���\�L�[�8=�r�} ���<X�מ����֓H#�k�)��!��76ߪ9��̽�׾��)���ڙ�������Zq�N1v�J-p���(��yu%;aɏظ�z�B
-���9�(��:lD��_�̦'������$�N�N]=-���`Sч�����������)�n|6�`�������i���|=��C�{�T�����a�-��[rߍ�K�̥v�8�}�\3�e�*ʫ��QU�Gk�-�ԆTb��A�_%��[��	L��r[�B��c�1ڗ�W�k��Ĕ��O8�/��.m���OK|��'�?�ᙃ�B=,{�k��g)�L&ް���ZS>�P39A�i�'�_rW�:`C��
ey�.�w��l�s)t=���o}N;t���AT0@
TK�9����ߛ�Qs(JO:����b5�E�V��O��Jپ��P�Y�v�>T@��n	<-7��8�����|����bo��}��|����=w�IFI[̖!�}$�r�~�� u|��N	�A�R��l~CI�F7�t`'ǻ���8P�`����">>�7^����QO{��p��`c���ZK���}1т��<m%�����M��MJ^H�Y/�[��/������c'��S�9��\}11a86����o�{��>��e�%�K L�|����Q�X}Qﳒ�i&~�(�Kg��36��X*���	gj��pb��|\��udוԡ#u�M�G<O�T��k�vw��v�u�==���3Dt���3%P��d�'��֪�I�}Z��3 	m���{�=��d�IQ{�R:� �"�7~Ԯ����&��T��E��c��|:*I�XI�RUϒ��h���w�ef�^^Ɛ*d}��KVUW���>ċ����T��; ��"���o=x9�dMN��J�����0	U�IV��C)����s�]�n'➰�da�!�>ٽB3�����M�Q�rǌ�UA�{�[��bM��3� h����J��Um�䩴��}i���_�,��nk�~w�D_�MQۓ�RlϦ1	��&Q�gY�f�|*��w��8J%���_�����D��p��!Q��8�Z������G���(�gA�Y���&��f��"�GPm���1��t ��)���&P����ФX����8�}�@?��}� Dn�C�����l�G0[�*�I�pu�'v`4�;6��b8A#,l�X���+}up!Z���Ы�ʰY;�O,��3�gVf�b'y���q�03O�ԠF�h�d�ܨ�,� B����ӫ����.u��F�z�agL��jb�A�u��zwͰ�aZ���23��,(3~l-*$.d�$i�@/���Gmt�<�!	�ɒ!�JYm4�?�:=�7�,�LN���)i%�/��i�ѵ���~�U_��\A�W�$]sr��Z��/Bx�?�'O��(Jr�ɫ��H��l�jykP����X�Z��x�\��d/;�1��#���)�,������ɸ�Y?$>s�#�=�>�"�~V��E�M����ۜ�.4���Z�E�T6.b�`�-�娹EF,��l�����q�C��-�9	CB4f�c�Ҝ���?x�z���ƨ'�B}ʲ+C�߿?�l��r��*1�[<��I)&p�NϿTe�3_�/�
2��N�����O� �b�-���4>����M#��=�s/�.�s�w^l�E��{Z�:*ĭ��6.L��T�0l �>b�K��I$_9��Q�)�����U^���Y%���L��N�|��B\?5d�c"�����B1��j�=fU�Ã�*5��ի��6s�s�,9LT�'���?5w���7Q>�X��+ �ǛQ���G�4wt��b���ҞU���]�zG� 1\��e���$������2a��T��+|դ�O=+���r�oaG�v��k�໶p�{�7����x�8���S�nn�Ƭ�r���;��{6F]߳Qu�b�� ��Gw�r�	j��v���
Q�)��T�ظ�A�W�i�	̟��i��Z��(^�ڮ����#���Z��w;]�v;��?��b7:��_�}��7z�����kٗX���g䱁5��Fiv1�,�w��b�#�\��@Ǖu�(��[O*&R7E������Z�����ߴ�pO?���r�n'k�J ��<���%��d�沰�ar����N�i�������\g+��;�������Ȏ&5��4�}�Ϲ����z@��+L�]���2�Rc��a��r]\�:����s#�-�L����Iޫ�Y�H+pD��ue�ǎ`k�uvƞ�''J��/yBwpUǬu5v����n�]����^�r���W�_�(�0����#�� @=�����-#�Ÿ��Ȗ{G��M��A {���j7
JBJ` ��������ϧ���VS���ލ��t��Q�-�����IR������;;����#���W,&І�TLJ�k�x�ka��6�}�h��]~/5���>)�񅜄_m���2�Y��K6�m=�B�q��w!=`w��f�_(���5�G�4���:�-H�&��i�?[vM_4�u��\����f�X�N�����ߠ����r������FjL�ve5\NI��ƨ�W�v�P���J�"�i����Y�i/��((�	\ʞIT�=���~�!W��ը����u� �Jҿ
�k��
mFZckDI� 2@�ܼ�������P��H�B�*��r�d�$���r�'ʴ�u(It3�n��Bc���R:#�q�m++�事�a.@�Ve���^��5W.��ޘ��i���wN;r�
*b����s��w-�픾q��y>�&U(��j=�+qU�3�.� \cH��Rz{|'��4����%/���g$Ӈ+ �:)��n����۔�k[hT�'���������-e��h3n{��Q3p��f~^L�%���R2s{~+��Z)��{t�N�qΩ�Wנ��|"[��+��m\��۫r��d�TK�+��w٪�����NM��~!�0Q�����̈́����v�k���`N���8�U�77���`��CR�E�VI�c�8U�F��lٛ��*&�����P|xF�}�F���-�@���:ʈ�»��-e`��6E95�!�'�m%�4A�Y�CU0���!�VX]�xA��a��9��~�̦Bl���u�����!M��!Eϝ;wS����L��( �^���/���q�`��̹��	���}?r�Buk��u�V�/!5~���8�x��눻��8��a�Omr�ӟUp���O���7,����m��u�4�����׭r��4&����M��OQ��+��>�	���$���$��ٔ��^�ڠe�u[?�ZaV�_A���8�D���sV���u���+)�zꔒ�ה��;aw��H��2R�bh�z�����Y�{"��$�$������ܔ��h"^|9}!Nl]��o��Z�͋�;�f�&�jd�`�¢��79���5�X%B��b���n�OP���V�v�0�An%�o�.�zGqY�T$d��E�U��#6����wx��IF6������~?M!&��a���T�ep�QT������Ī���D����1�= @����u�;l��ZIM-�5�@oc���� ��~t�ؗ�nN���(��`�:9�y� ����ǧ���;�3�3���C�U$���;��N�p�@]$�<d�\(�vm�,@��ͻ:Vi�-���,aX�����EL�_�[���zbV�B\�C��&.铼R��u)�9�C�?~��X'{�q��)�oF"�~4�KX���c:�@XĶnd<����弭ٵ��ڒn���{.
��)e����,�� +N���y��@�-��HZ�[�s���U��Z����~��ߺ������BClTz@��;�G����&))�Y�����=��]�����ǈL&��c+��#m����V�Z�������R�#����'��߯�{�Aՠ���4�N�68�[k�^Q���\�(Jmi��Z����U/<J����{�f]21گ�N�Pm��c�X&�R����77/d�U3#q����E632�w�g�
�aA��xe+�zj�0di;��ǀ�ѷ�ځ���J2=��xd���ލ�oX|����.��q��%N(���/¬���(��f��$(�p����WjR�V�X'=�}�70ISBL�M��){���{�[nK��x��ݔܷ�HSjkj~sW�zzspk����82�<�9vq����}mPP�l�3���o���-$I �1������^[����E	`��b5�J� 78�#!~�4�p��pp�M�[�҈I�i���������:�Qe���J��9�9������ǎ��FSn�,����$ѬfЏ�X�-̈́��%7�^����K���i����y�ט7�ufϟs
7iv@|)���F'�&y���+fU_��?��VZ)͂�:9�dBH�,S�\7ϒo��e�}�T��i�ݓ���\��}Q�=�ym3���T�0�Pj��g?ͅoqL\�֥��<��'��nʙ�eݭ��QW�'�5p��Yt����y�6Z �Ju�-����@3��xC�Ԇg7�&��8�\L���/F]7��"=4FO�v����_'7�vB7G��k���GmYo+��p�g]3��ch�� 4�4e���̦����ʵ��~�2�,��h�0�/�s�j�w�4?	4��3;"TB���B�����
�qB��r]��y���$�t}"1�R�
���On���\�WP�'NܭW}|���0��s����N ���DtLQ�_�w1��?� ��>ߓF3�L�h��쮡;���n2f%q
��������ٚA����̫��cB��;~�{�]��)�ØR��� �� �6W�,�m�z{�,HQ�Y�̭�XwD�_{b�F74f�M��YV~��Ԫ��#+B�6*�zB&v��6�K"}Ǫ��E����D�:9�8�� fM��Q���Y���M-H�%�%33�l���a��K�t��r\op�����uz�,%)�S�\mq��#�݆���V~�V�)&�k.��������n&�z��0[%pl�H�[emm(��ז�N&G����a-T�mΏ�|	��w�s�!Ҿ-S��,ec���2Ǭ�-C����:G����@U�6���-7!	�-[V�<�w�:�3��\�T�΃�*(_�w;���--��$��ގRu���o>\?�ag�HI�Q ��#���S��G�M��`v����l�^�1�;���+�PW-rbp�Q�￱=�_���_LO��5iJ|gU�%n�	Ȕ�z<�V����raG�}��vyB�v��C|��5��N�22o��$y�jP�U}�rJg���来�J���y�؈����W�������q�v�}i�Oʂ�hcko1?J��l2'�+�
Wf_ׇk��/{$s�o��1�'���U��/����ˎ��ʬy&X���r&0�`�d���Z1�u^fmZV���VR4d4PO$�����] 7�)?ғl�"X�ӓA���<o��>[/sL̑��"Ĝm����_ژ�q�v5��VQ ��M�pn���,M�M�91h�����9�N�jj�P���m5;.�<Wb���%0u������E_���k}�֑C�M�G_F��ɘ��T���JA�.��3ZQ�����1�b[-�ϟ�Bf�vgZ]�Lks�+j3U�4���Ri��p�LLH\�=�#�K���e,�W�`#n���`�ڷY}�ĳ�~�It�G4��^s&~��$��ʢ�1kI�5m�] ���Io�뫙M�"	��:;�43�T��{tp�<�^]�rę�H���HV~����v��w-��:�W�Э�j��� ��v����\�t�ɢ�_��fHE�]�@wg�:ͻ�&")&}g�r<��ت���Ù�)ٛ�gc��4�N=��!����δ�m�LH������=U�$z��d�V9�n&ՠA��9���fZLz�֚U�������� ��q�lP?xBBLLLXS(w]i��x��1� ���?Ko6?�� �k�<%i��g�M���Z��PM��6w?����P]A9��rOT��h���6��[��?�9X�C�ķ#Vs@[[���鿨0�ٶ�7[�h��J��mv���ĭ��<�e�;;<���������-���_�b�t�J�8I�IR�y6�M�k��Մ���#ް��[�q������Q0���aݝeA���o6�G�z?.�o߾����oK���w1#gt����@���p�\���PXGmJ��TGQ���w�lo�Z�ȬUVV���_������AU_D;��L���'�4�^�mN!�q5��W�V�By5{��Qu3��?���;�W��aI��kս�֑2;"�W���}P������� �Dc`i��3/�����<�|VP���W�K\�R8EΗ���A�mKxۏm����3�	�x���L%��z��dM��sw�V���|΀0�]��[\1~���φ�W���g��2QƎ��XXZ:p�D����%$\�z��?�4[&g�xT�??���x�K�������1\��e��A�޸,�͏2A6ZS�2O䳾@��������w�諭!aV,z�,��a�󰺯/��E_?X��U=��rخf�eE��cZɝ��^�����&�u�N�f�V�?����(Z�f+�5}&�%���0�����J������r�C]�5E]�(<�\_�*fH�F��RsG�K�Uee;�����y��d��^7j,Qz��Da�l�o���W��l'{�z�c����5��γV��j�����~X�����~*[����@���C��0�C*��-gs�ۡI	��[���W'y��%kM�h &��o=��S��QT�z�k��ͻT�5�����j�5Jw�<��j�ݰ1���?�j��7m�^cI���柶���>��ӛ�����`2���WV����h�0�JP^���v50�=�W�,
�i�u�2ϊn���Y_͡4��g����ޝg5�����J�F�ƞ��Ih-wU`�[��@�������~q������q�4�ѠYv�F�`:z�=ڶ���m/rtt/����,^��-GSk^����}`#cVyT����A���cfG���k 1��,��h�� Ć���sT��^7�n"-�[[[ۚ�P�[u~�\��Q���r��34wK9�w(�&ǥ7[Q��qw��pvMO�Wbt�r������Փ#ீ͢����Y/�UZ�ڼ��j/m�IW���_�zx�]�m�V韓���ыN�{Yt�����g��"����� @���%�w�7G�eoJKKF���]��ʇ�n���(7���L���h���C^7�L��z���!��?�Dv4&���<4M�f1�O���L������\���kw����*/�K ��Ä�@��Q�<f�ƙX�,��_�������oIМ�3Z7!�\H��8�t��c��ٵ� H5���ɡ��)��"m��r+^�����DW��������K%e�dc�v��e�����3px�փ�F{�|���5�ZU�}�d@K�$���R@_���k;�Z�R����(̖�3ت����z���3�-������c��(���Z�'<���{(҇͢!C��(�`v=<r�wrׁg]TA��a�Eɰ{���p�q�(�$��6� g�� �(������Ҋ`ݙ(^��Ue0S�dӶ��j�1�8_�r9b<؅!Z��E�Y}H���"����N
�V1���c�A��!� �.]��W�� Ǭo��D�r&]!��s�Rk�G�m���PK;bӒ��yg'�����1�����J�QР#�������5UG�"L3׏�t�����c���6��=�S��x�f��u�����Ց�U��C�4 ����U�|��*�mE����L����:F-xFF)>1����vXтE��J^7����9h���ş�Z����^�!U�� mΩŊ���5���ɥ$��D�Ю�c�{�JwJ��Mt���foB����I����%�mmQ&�eh�e��% ��O.m�2�����[�j�[h��O�~�B\������s��#�0��?���XCC��xs�5�������%t2�m��.���t���\�%�3�dPe��oh�{{�QZ}��w#�9��}�I+v;'��h2���u'x�8�ë�OOLP��g��-�4�鏺�==)��yO��QK��Oe"�L�t����1W޷m:0W��1k�#��/���w|�P�M����[wjで��t]���@&����|˻��[�n ���	D���U��~���5�ݯ��|)9y݆��D�AwS�2k��N�x���ߡ��z��]7	
:tE�N���Z�����/��x4���\�����	���H/"����k��=w�G�1݂=�=�]�W�*�"\��n�@W��r��G��|>cC�U���؁�A��z�%RL6�#���Sؖ�Η�7����FQ�IC�QO�B�?6�R1�����<0����l���2�q=q]�e@B��ܪ��lP{�l����ߚ�P��a䮙_c҅{����ʢzO/�w��i��<7��uo���Ǡ[���[��������m0h���C�ʶt�-�'�=6g4�R��>�j���O��a�np��j�%s�l��s=���(�%��w��/�����K�E��U�j��;��!S��j�U)~xPNa�׺os_�}/�<Gȏ�ߩ4�m�##�qܼ�-�sNU��k���$\m�i&.z��4 �3��i�elKf1��[Y�1:����'^�8s0�K_����=����ׁj1{Z�yn�?^��������^ءk = �~p�1
[ct^�C�<!�s�M�m��	���u%M�F�V�Ȝw_
*5%�jqU�?�G=h�eU�����ʟ=��)
��<B��">�hhG5�d`L��g{����F�t�s�&�����@׋Au2��=�I)����1E�>�S��EA���zu4%'��U��[��;��Q��y"��.����cN{����L��]5g5��lʴ�s:���R�`�XJ1,j}��8�:N_t(M}\�=�EMI,�m�L�)����}z��H��6��Z�ͩ��g���	�
5��*���?m�����ϦR�ZCc�sZ�b�Z����k��P�Px���Z�Mh�gN�-7H��$��_\���}���.����ɩ3��[�배��0_̌l2��մ�öuS$\��;T�� �wv�.�%T�S�i4zΚ8�}�>���/���� ���,�\t������>Y�1Êum��TVA��=��u�P	͵`��M4n�cֽ�.d�T��*�W'�#�?|[�ڕ��:u@=�@f�r�����3k���ٛ�j�|vd�W'��R���dťs���q�mT����R�l<3Q��6��F���������74d���F+}봒fP�1��g�Ǳck�ПȎ���3��e;آ�3�h_������Ϻ�ﶝo��j�#�O�U-0{����m����xl}K�KP�P(/�W��T��J����E� R���Ë�>���;���ԬK�뛛��ҠN�3�c姕m5��k��zs#O�J��	 ɚ���l�nn�T)�&f���䶝�����w���;�d�=1�2έ?���C�Y�h�1��hO@�R|(�בت�8&���*I��hAy��d͜�lt5^�����&�-F�������Tj�1k����#�5s�!Q���􎚟x��5G�A�]>���!%%e#��ĕ[�u*'��ɖ*_�Q��U$Я�x�9SuZ	��vu^l��D@h�w���2��C̱�0��W��<�#O��2��ܗ���R{7^��,�9h�l�B��t1hL�*��9d]��Y� .�?����)�JF�?}��v�ً��lm��w)��S~�	�+ٰ,Xx�K���`XJ�kP���c }-��Unl.�/���./C�-��8@\nQ�*����v��W�U
�i��ϵ����bΈS��l��q?<�,޳1j���H����U���k?�!qB��b6{�=2Q��Y���>������S5�U���B���i��ʬ�ި��y�FaY�(��*��Y����rg	/6�a娿�!��9�xrB%�]��(�j_k%��T�IV�B�}�N ��(���pi�^}�~%P���K�ǚF�z�/��K�y�{����uuƯO�^jgn ������a�r��M�:�u?�������uzӢi�,����=��W�iƄs6��j�Z��6r+5�̳J�٫�D�$;˯+Zˋ�/y���bC�~�,�uoX�����ϋ5L�D��ۼ����f8q�J$M�{�����=}�|د���.�8����86cO���Ikߜ.�r�#���J�2j��7:��Y-��/A��N6�1,�2���ǼE���ѿ��(s$`GVys���C�75ChdA#\��ٺbAP�j�fwf���H
4?�,�ׄ���mUT���a�
������&ܮ�۵���'���J�i�Sb��P��#��� ��W~��v	h�M�Ú���?߂����B�`/���h�Ώҵ�����je����"�%�5��bw�>+���>���亊��1`����t�� ��W~K�6wfz(s���W�|�4��\�8�0{SY������y؎��U� (��Z^O�`[���(�`[�ǉw��ʭ���^�l��z�d칾g��x�M�U��6X|^�u�Y���ٍ�g�e�S}�?�T�^�#�c�W��2&�W1�jB�`���~[����� 7�����%�k��h��X-F���ޒ_�ǳ�H�-��`a�/�/�T�e8���M1117�yB����<Y��'i���+��uק�Ŏ�v���H���z+u�E ���#`ki>p��}b�g�܄^�Q6.B��Oɬ��J7)H|���>���JژE��܋�������t���Q\oa���P�B�`�=����A��(��F�L\ܪ�=sq��4e�u���γ�-���P��pz9ۮ��,*���g�Ǣ��;�sq�ҹH���u���i#��O�L�����m�z)&��rMGG��n�Lo���k���PH^_i�k�����ZN�I$�åR3�.���#'�w��n�wkPf�iP-�����a�xݴ�p_��{'pe�����,��TU~����V����@LB>MC\�ʎ��Q�ڣ�zƞ_G��SB�	M'|yἼI���"��ǟZ;�&xl�� �^���鹮�q
GQ�~�[׵_���k��
�(���b�D�*7��D�#����zPl��xѸ��P<F
$b||��-;d�W�P@��8`���LkZ�r�0���.��g����6��ݢ��^� 2$����"r��L�rڐ�TL���%J-x�7�By�hdw\i5����%��U=׭r����Dh������}�ө��8�=��=U)d9�CM1G��OU"Ӳ�*B||7D���}am�]^e��Ǳ�<<<ĎYS�j�ȁ���3h�ˢ����5������K�"�����������`��s�:�m��u���2�;���y���VKkk�r�@8S*8r���|�o���$/�@ؔS�Aa=���o���8+�E�d<����8n15������;:�>�j�yb)62�6��� �G�n{��ޞ�������v��8e�x�.�4����r�F�![斖
�_����VA$kw�S]�5����dpp���ڤ�s��Z_�{6��R�P-�r7����2mq�Ϯfp �0ꩤ~�y�IF7�sP�R��9G�'(����A~�Ip�6�m$#��p9��nE���μ�z�#�_M������G�	_���444��co\P���r=�v��9�al��/�����W>⃔D/�~Iyr.c��9�K�0��[���6�ܒ��u����wx�������B�>>
�H�[V�h��Ũ?�wiJk\2�u,�#�#��΋���q�:[���^y|�Ўޑ�4����J�'�0Мg?4PD�3�*~巪��uG+��c��|		�nnzj��}��?��Ah��!r�A��"�f�ةw)^�W|)��٣TO{�w��v^���ȑS���$R�32� �\2e���|���uoI�2����'�gtGV��z+B��yg쉞��c�*v-Xe��(��(���M�+�Q��@�DP�n�t�X(����R쨈�4�&KUpi˲*"T��Ez�Uʮ�o΃io���}�$	�y���}�3s���7�}�A�i�dD�-�s��� 狳�C}�����L,��}O�5��5��X�ZU��~w�{碘)�����`���Ud��Tψ8�0�� �ϟ/_�֟F���Y��9�֚��;�����-�|2���~Q|�"_��\���z���!�	��Wj6�S�2׬rG��]_f2i���&:{�8yYv�C��t~.A��6?S3�:~whpv�O)�Fi>J��P2�������7O�H���	��ϟ�k�~��Η)Sβ��z��֒�=�>�`�A:藉�S�^���Yתy�����{m���u�Cg~�'~�	�y^it�n�͒O�	=񴍌�xW�d-x�6�[�0�VM	^=_�Bd�ul����޶m��\��a̯A�x����0���-q�(SwY��*G��>�&�v�.�q�GA��ݽ{��*��Fs�}�?(�ӕ�f�s�h��v1�l����؃H$3ٛK|������h���m��&��f�v�����s�R��G)$ZKQ#W�.� �:�p��t���e��k�y�J�
�U����X��R��:�+ϙ�GT>)�Q��ӿ[|N��cn"�'X[1o��� 0�Q��/��,Ov\�A"�i���P#^�����������±��KEh�*�B���ZXr�ox���3��ۑ1q�{3�]�P���κ��5Uy$�zJ��wA��zXej-q�� a���Z_ ;^���S��/���1G�a��ZX6:�.u K끟�=i9�S)�ߚ�kAt���653C���ǨLb{� V��!F��������`l��7��CB� ��W�}�����dAHE�b!d$mG�M�=��ޜ&��
�9����y��~-q7��7�x�e�Y̍J��ow&� �x���E�<��Nɋ������{ "�>��[���\�6lاiA�����$��Gư��0��$Mq�y�ن�_r�<#I���h4��./�0u�S���]l�7���&1���$G{�[n�:����������&Q�)�C\&�F<N	�_|6��Ϯ���U�����uw��L��~;w�/�쌃A<�8�]$���Ab������V�-*����xʎ0+��fp�ځR7Y��U�ܫ� ��x��>¸K?��'�)>P���3��7ۈ����g}/�~��՗�����y�Z�#p��s&J��PJ&���GW��N�(|;�n�����OT�2��Qt>v쉗	��c�W���A�}J�9���1{ɈRG߱��p޲�An�8�<�q~�#c6���?�!��sȱ����ɁTn���ݴ41�p`�@���+l�d���"3b�(����x ���w��V�(x��i<'��r�����!��W ��MPf:y�rhG��	;���\tN	��w��m����������F���:6�2�DJ���D�}FF�����v�W���HT�N$�Z1�j�,~�l߁�DT�!�Y<S�X�.j@��W�$·bps�rr����>��h��/��#c?�A�}�kW�y����N�}�(:?�4�9�Ls6��@��ť���=hZe���z �#q[Qɇ���޼9�üP��ƶ���,������i��4�R����PLۑ��E6��H�l��zt�2c~J8��zܡ7(��(�(Mg)3�0�y+2�~��]�l���!Ga>��i<g���ts8�
�n"tsm���*��_�3�B�חѐ.��Lͷ�B|��stSe��q`���L�>�zڎ ���M�e ���<�>5[�=�^Bސ�8s���fY&#�����>'�$r

��f�bm�öl�r"�IOaɚ�CC�M ަ
��e�@y`�a����c#��$�^,�GB:�w�[$������D��k[�ր��ɾ��5��K�Ø�e�t)��0��h)���9?��f�+j�B�~�����zn�yaT���!�R��	/���T���r7����~ ��
�CD��'�⭴�>?	G�7��Tt�]⒫�g�JҎ�2�ގ����\�����HFV��뛥�����d�ռǧ�wkطW�
>�gz��?twp[e���%��S��2:<���/��/|�[�.�����>w�Y}�pW������qs/dp�FY���'̜e{h����7BdY���,o��R�t���!{V��淥��!�����5��AQ���+��z�[��_?�/)��ie�5�;��c��Z�Æ��k	��W�9S��=���F�C�T(��!C6��� C^��y���Hj����W�.�xD� b>9	}:)z�ݷ��'
!w��܉7���"����P��y����&
���^�AL��L�m 1���NBE4�F ����y��Դ�Ɨ#囹���ؘ���"䱅��_�j�!yH�FG?H9Y�)�d��r�-�0 hF��F����uH	�&`������_*��>������Y�6��Y>ɜ�s�����i����AnG��uCX�V��:�m_�"賣��o4�o:'f^Gr[ݣ�Dt��Y㰛v�D��)�  ,x�^J=�����o��/1�,e�����YDژr�Ύ�ju���O}�fۃ}�K`�?�ط���Λ��h
.�m��8;�
�����h�"g��iS76@	f0K�Q���J��`8"��c~��i�e�O�����F��'~^�zQph�B��۱�΋,�[�}ʖ�Sq!2~���;|��L!�K��,��d�;m����z����`?ﯟ�Gy�?�Nd��,l��ze1ˤ��B��8����Ծ�]��(��ݧ��E,�/`dv�{��n�m�V=�L�n.;o�_��З��|��N �~	�86*��{\fU��䀶���\��� ���#�A~?c�k�-t�;�}��Q7D���ϙ$6Q~`9_8�����lh%���;��x ���<�0�]2&:ӕ���_�>��&�	��(�K#�����w����R��o��/�%� �M��u��Q�	�������j�\�K��!�Ͽ�0a��R/��A��w�oR]C͸�/%��m-"`3����A�s�:E�`T���HA�;P������ϔ�܄ż�\���q0��Xx�v��0ǎ»OgQ�Y�?Ⱦ
���񼿛��KX�7��~�:�3QH���"OW(�7�h<�X�ψ'w	�=��M�Y���Ҧ��"�rt�|Ş��̅�x�S6���1Q�����F!@@Q˕n�����1���؅��NՑ޿�3`��z<�����B����yǼ�N���s�6j���k����"~�	d�L���$P�s��$,���[<h @�99m��d����䴝��VJ�Tu�@��߳ʟ�s��t���e���<�<�=�{c@����`Zx�:YRR2;s̮�}<"�0�T��E!�ζ�r��*���A>Y�g��6)7�^�������\�_*w�Z�!�b F�fVȪ���D�7QkN�նHÿ�&���� ?vѽ�8uS:	��'����@�&[�K����:�����Z�����E�c�]=����CQ�;��ѽ�!�'�M���n'�&�o��>�<!���<VV��}�ӱZ���_Wܥx掽���Zٌ���=w�m�m{#&�k*���?�����f;��b'R��v��D
,ԩ�'�����>�
9�=�))-�q7�}X'�.}����;q�R��A�M+�>��!c�:�ԥ)RRwRH%R+ɜ�gT��;׏�]�#�g��J�Ƿ�����Lx��-��{�l�=��u�b�y��̳���v���' �Z*X��mi�'N���N�{�|oDdd � ���Ű�����E����W���\���^���RU`���!�qu�fZ�W�c�:E��-<ɦ͋.�f������3���f$__E����$ny;����vLHR����U����q��Z�ҡxO�٩V:3S��spuu�t��3��7���hQ�p��Gl��7O=g�I+J���o�X2Ӱ22���ә��T�cb�嶕���m�vW�g��f��;�įJ����.�Z���;0����ć���?F���Z���Y�8�~S��V��MRٯ{��f*�u`�͖��=~ZѾ��>�.`�M@`��A���.7�s����DdIg���h�@%���<��a���D��l,_�7�&��aK�T�c��A�~o����K�ƥ��;b;Q]�4�|f�G��4�F�������"�^��&�o��ns�=�(q��׻�m$!���F�ZR��f\��uVD���O�>5��| ��k&�0�q��w�
M�h}�;d��(��8� ?Z�/��2������h�U�nF7��3-oq9C
����x��M��맼,����_��ZS��ͪ����E���4�q~��:�儨CO��f+KUGޏ��z5��1'R$m��{3H�����V7>%�ˋ�k��)�>�����b�1GL9�=�9�<���uH�w�jY'U~�N�z��j��&����b�cS~�e�#_$�V������5�C��xH�X�5��U��{y�.!(f���6MU]O���e�#�p/��1iDv�Q���{F�;�;�U-++5�~���$!ǁ�fI9��z"��:	��(��O�&�������?6�\԰?�d��K=|\�-B�����=.^Jw��&mɶ��t
�jP���sl�QW�d�Ƶ��e+kٛ��9_��o˲|�O��oN)�����[���7@�RR��=}|�Y�3�v��CX:N�:FaO��؝��<׭ł8�=_�tӼD����'�!K����]~�RA�۷o/dH��U�i����7kK�u���ÿ�0�ۭ<;��_�L�p)-U"׆R�x}p:���q]�M�(�Г:�����_�Y���_C����o��j��J*z2�-�D�`QqqB���c�_In�!�P�����x�k=,��*k���^˳g;�R��9��OzE�SN������O�!��̈́!�d��_�ݽ"�6Bo��\��
 �̄1'ߴK��D��$d��3�%�j�l��]i{X'K���n�#����Y�ý8�9�0�L�]�;$2��a���&?�(Z/���)�\��	��x��V�����US��e�6EA3S �%�b����r]:�>�
Ǔ��}����ȫ'	��zBs�����r��4��g��1����g�����V-���*�w##"�Sm�g�B�ibƙ�H�||}�w		�O
���W����
`	�K��z� �Y}$�N@)�Wmd�$�1�!�b�������gC�]��Pt� �w��[������������[@��U�|��4���s��y��Q�r?�K�}��kך�~\$�hmê�1Ww�7���z"|�L`hg�5~"�{�B���Ǒ�)�Wey�^1p�|�״Ml3���:6��t�<`vJ%f�N�_�,Ñ�:c��Jy������QC9���`?�o�Q.�����t�`�����7�5U����n�3$$dX<8H�9�������L"�oH�_A(�'�gF�ݏ�����6�Ē���Dq�<;[�H33+�vS|����%l���g}:XH�n��Y��G<���',��B����S��:�Y�U<���rT�Q�����n�t@�ɷ]X�	�&u�V�����B�{bUq�q��Rx:r�+�����N����[g�.[��u+�=�~�����˯��N-����?N>�uɗbZ���dީ����,�g������Kj��Ξ���@��z9��Z��|�]�~�[�'KS�\Π��_�J�=C�2IK���7U{~q֊�w�,.*��zOq���*	�DIl;$���h9���p�I�+�[������qP��lZ�=8xyO��A�$���/y�ͪ=ɺ�G�Ů�ȇM�w�Q¹�6ݡUc�����N!{�:Q���p�,:��G9��S.9BD#����}I�!Ok%�a;X:Dֵ�N��6�˧�B��s��=�4���r��]k�i��wM>|g�L�P^c�l��\�����p8GiC���O+t�M]����@n���fGg����n\Z������������P��AC���p����F�??{=�TN5k{'��6��ZYZv?��!g�7�:)\����A��}NK�g[ϝ;�Xu��`�衜P�������H2TU�+~�����7'_��D#v��Wզ���,����f��j�,s��g�#\9c��z���Mo��]ᛔ��v�UM�g���kש��dF��Q����j�8��HD�G��\��qQ��N0<hb� jk�q����ϊө�yq�һMM�k�'e�y���ͱ�M^��jG�#��o���خ�p}������S5�M+�׵�i����3: �`H�Ό���<�
а>ʉN3F���I�d�7��$tw�p��(O�w�j�ԙ7!�\ѳvO�P�
��|�9�+����bD�O��"��x�\c�0'�lm���ֶ�ef�P��=z��	��d�t��������{�"fS��0�����D2�l�(���<ݰ��^8[��o�݈�Q�)G��9�\/54���$�t���MH�_��p����X�k5?7�9��ޜv/u������8���jY�J~A�p�p�	�A�&@C+��I ��aj�:fҧϳ;���H�������
E�v�}KJ[
��z	��v���>�@D���k`�q�u�� H���g*٫p.�V_5x���UZ�f�im�,xc������}�F�.���M�����<��I���[�(��6u�I }5�-l��t���
�Fi��{n,V�(a�#,h`�Kb@ޤ�������o![�ʾHM�ߒ���uH���a^����~]��qJ����u��Ō��D&|@?���fWX����a��6p/����Wd���bZ�Mu)!�-K��g�ƍ�_����Z��틍�Ǐ�ne��O���ڿ�Ɠf*́u��������L��|#�#�q�-HI�yP���)2^u`�XeH���m�|+�i�!%
�n���T�@�N�tx��g��������m�r�j��]��D	�!��D��e�[N ����� �I��_,�o~�@�kO���m(~�=��df!��fp�^*�����~��5�:Ғ��9�Ϝym������S��>mr��{R.�� O���1UsO�o���Le�z�(d�������LQ0O�]��_1�ͥm`�@X3]8Ba�����V� �~�}� ��#��r�����Ć�T�vIII��WWU�:iw��=�?}�bff"�|�Y�(l��,"�d��2sBˉ��JPIR��� ,�˓YX
lXF��m$1�f���Roy�|)�k/L%m8�;�O�{����{�]S?]���ԟ|��9D������^��HU�R.ٱիl9ZYM��I���ؘ���ؚ^�&i��&Y��/�锑Qnb��)
�xc�RVSHqq�3�����y�+`��_���Rh��Hf߈���_L����L��!������nH�d4������=~�'�`�mc:��ئ�@H�3�| �4��.PM�{A0}˥����U����P�z���Zq�w$�qG=I<�s��TQn>qF��$�6#���&�ފ�Wm����4�L���w^[�O��.�u�������v1D��_["�D�.-=�Ѫ�Tz�UEz���B�v˦Zd(��GVf�8�������,آ�X��Hh�!�^��
�U���Rj��%�C@AR����9�J�<i��);�	���\�@_�go����l��J��Р8��|R����V8��4������iŕr�������!/�����}
`O��܌����a�d�4�O{�����Mot��A����FE�79��ș��K�>�Ў��QxM��Kv4�Q�8\Bͧ"ϣ[p�e~��F{��]P�����V��6���䓉�\����<)�챮&J���������j#�����*�Wt=�Y�.y[�����i�]y�Q���D˺��[����b᱑��!;�H�F� o���|t��3ajxO�r;�v�W��u���s_�i d����XYMu������>�����E��x�)�;�#�]}bC�u���{��a,�v���_��/)�R�*��C��w�'i9k����hs�b�ľ��-V4Wx�Fu��/�T@"��W����G�l_�\S��x�=t�k'B%�ܹs����+a�E�������:�Έ���tiY �hQ̖��x5�	��C��+�ۿT�<��r������#���4
��]f��׵�9E|//��)�R 5��?�PMBQ�JԌ�@�)�:�pԺv{ooS�+z=AU1�1�I=Lm����2��X�(س��SS�� �c���u�� ��5+��Z����*�����'^���Y ���a"kG+�N�i)w�.���"EnIl�zT��P#wjP�"e�F��Ҽ��������g�̪�+��dN�g�0U�F�a��
@N����zl�H����A�?�x?X�t̀Ɠ����uP�B�n��$�Gc�b�hh�����qc(��!H��7@��œ� �]�5cJ�?|��H�(�eL��D+��d�i���h?,� R�n�hH;�
E�qu���de��� w*�����xһ|�Q��%` ���u
ڋ�[�=EL�{�T0�=Hb�,irȡ�竓?�3�])����)��3~��f�N�a�F��������@YYyjN���oH����轾�P/�����ӯ���[�J���5Ω'\����Ɲ̝�
�|�ν���ͯ�h�Y���m0�6�'P���}V�yt�Q���O'd���:���xJ�)�Pw3�Mq�Eė�B�A�8Q�65���ߔ�TH��I�bf�:BT��?o:�LC�)/Qq�r�XK ]�D⤦Z0ڱl!�\ĕ�P⎼��A�Tog��qS�����Cz��'�Ĭt�(ܢ��:һ,��A��Q��UG���Vt�]���+Z9���c���$]��ܽK�5	}�'f��52v
2�I@�]wM^��z4�C�t��[+f�}+���+�; Og&�Ls�.w�jҺ��A#	�vR�`/��	����o��(�~'�D�A���{A�Ǒ�X �'�(6U�0�}Y}�
g�?�U��xZu�9����N9qu,��>ĵV��p�v�r��^����N�?���Ӯ}��B=.M����Fu��T�/�1F���>����%P
��p���l<-�U;�h�/��i�[�xZ[�5H3�²�}���t���M�M�2@/)*�����(O��ڍ�������5���c��+k��G�+�D��}4 p	T���nwP����N�#��#�~	h瘝X9�H��u��'�q��-P�
=���g�G��6m��񶮸�z���Q��=ޚ3e��.�0ߧ ��V���i+�e;����6F�m��}�jq'�2��"�N����;�Oۂ�$��{���3� W!(<���QW�eL1�)
���t(�"\"R vA#���w}p���錱�i]�q�������Ԓ9��¥�|V���dN��`����^1�a�������,&L*��i�R�j[�D�GMȇ���g��(6���D�u>����\�Xn��xB];��2�X/��׸zO�N���Z��&��ߩ	���{c��lܒ�6[?�7Q94.�z���6�p i�o�siާ��XH����&F������8��!�RǍ}n�v*�HvC�d������&�(�^�LY���G�k �z�-J�Hk3A.^O/�=�G�zf���,F���g]��d��ƼL�Y8����K �����i9I����H�۷�j����(�$s.�&�tφ���%3����}A�q��vRx<�(�^x`Q��������:CX��é[����i6���y�<Iu4��m[!_h#�?�T�#ŝ�)�,~5�h�p]7�' �>B.�������j�}�8U��Y�_k��٤6g��)����`^�X;`�ӏ��p�����a�"TRߞ����k��`�#a�|
���4��٤�F��F��Z�����ņ�7+\����v70K�IZX���υ�9�2�o��k�Cn��ta\ �����	A�]8J"�O��du�T�숭�Noq��ڙ�ZZ7��=��ˍ��]LK�@��(1*q3�*'l�lsZ�m�z"��7�n6�yce�
�azc}��"��#�=�<7��ɉ�lt�Tg~��­W�/����v�.���M?�P<����
(�:>4qXѵ�؉w0�8�� ��v�k��r�c���C�㓕ݙ��E�MƢ��!�	�ؚ͓9B��GoL]�I3��Yz{���J^5�c�'��C�нP�'d�6�������5��=�V����������Gڃ����������rmi/�}�F�Ϟ*��ثY�s�����4 �V�ZU\>h�ј1��&�V^	�?>l���9�F����g�|)Dx/(s�u��ux���*&о�lݘ��p�}�ܪ�js	���YX-��E���t��]��{�P��s!��s5F���4Ga�%�G?�N�I�m����+����(%P �^0�*��*�	ִ�J���ДU��N��N݌Fr=��Q4)�:㎪�����Ik�-���=e����;�4 ��ѣG��Q�߹���[�K�Kp���]z��l��Ox���s��m�a�ӳ?D�����X�a�<�r8�����=-��Y����oiT�_t��d$&H��T���M��q�f��M�?����G���&��f�T�g+<�ؚՊ�ᒢ��VR��Ab��5�juڔj�Զ�����������u�_]���<tO��3���������	��fmC�>����x��pmX���ſ�uʤܯЪȜg[�㺺����I�hǋ��7�����m@P�oB$��blNbV\�,YO����x�M������/�~'5�9X�B'��5H![��5ʥ�	���2�@c�| �k���-n^ �FZaywsc�ՙ,�܃R�
����W���5H��P�ya�j�NP��ߗ�!*��
i��o���,�bep��n�a��M��]5��u�zR�X5RR/�$k���;::��׌򍈔�������ʡώ{q�����x��0�9�?pͱ�#�x��%�@=�ƜP���1  ������N��./J[ V�S�T3_]]�;w�%kv��݁5�o� R��_����q��[k�ǟ
�A}��D�����n�G�g�Fx��A����+$���J	ɏx/�K�P5��'S/E�6ިg��B�<�:B�F#�4y�D�pF��N��u/�-.(%{�Ī���`=�Kņ�����z�U�RZG�@#T��{��P{	k��$>(��b�������G�E�h���\�qA�6�q0Zp�U��R�DU�o����@�N�0l����y�ѱe��c�>���x�Q�pX~b�:�/d(ti����4�6������7�z�6�UYge��UVK�,3�ak	w����b��<��p��n�J�S
�����0���ꉄNMy�#s|c����7�����K~�����y���1�i�"OR7�F97����m�%�ki����>����4�B��}���b�f'���Du�@�n��I�uX����mJ�:��͙D��-;1=��b!�Ju��|ݑg���l}���v���)���� �dq[���0]�|w�8��0����!]��'i�L$�>z
�Pu4����Uh;K3ﱼ>�ŵM�ܻ�u�ӻ��x�Id�*��no��������Q;G���3���qa\��MB�1�n�6��٢R��ǒ���A��Hg0u��Ej
Ša��>��D�ȏ��5�644��Wԙ�3>e��|)ɵ��u`$�plOi�=��(Jp�t`��/]%�Ag��b}A,�o8���W��o߾�$ʑ�}y��
��ښ��ׯt�y�ǆ$�ێ���}�i=�Ap�;ǁq���������A��u�Y��էjC�2�Y��hf��#w��s�V|�O�1'>;�9#���x�W))M��~�@�J<�o��Q��S����Pq�u֤��^!Qz}�F�囦�B�<ߩ�&���F
�ʹ���f�8`���};��>�X�{2N�+�y�+���%���� �������BW|�*RI����z-��{���<ٖ�:+��yh��	�����CW{_��Ǉ�#ׁ�:Rϕ�-���3�7��U�F@Vn�'�Of��ͫ?)���ƀ�D���16a��(MZ�0�^��?b�0I��[��:�c9��n*)0(ȶ\v /zP��K]m���,KJEy��W��a�,�����͵V��U�/���'(�=�I�FmU���������Q�փ�E����̉��^1"��t9��J�ͮ��v�r!�UwƜC��f��R{��)���VEʑ��۔��jP�Z�s4!Jɯ}�g��Ϭ���^�]�v��rK�>$��*Z(7�D���ǈ��z}�����n�����,"�61����=3����f����λ��#$!)�?�G��%.۶�k�w?+ȕ�<���f&ݓ?��Q.�%�z8�m^08ȭ9��)=˲���T��,�6�M�k��g���9��_NV�����Zu����Q�ޥ�9T��h�Ag�ڑZ�r'(H]16��i��K}�%2 �p�#Ǆr]�1����yԲ7��Y����Z��k�~�6����
I)�f.	B�~]T�)�f�r�~�����̞���-��L���������ۻ c[.w�un��@l17�EV�!�ꜹ0DzWCmdn�G؟��sZ*1U$<i>B�ocQ��=ۭ��o�P���s���P��&���x��G�]MEE ��RMB�=��n�d� ���2�^>yuЮ_���1�+D���;�5NJ�Xq2����O����c�W���0�i���cYYZ��" � ��ۆԽ�3A��L3��x�-�Z��^BM�D|���=�ĒgJKo��T�-�}�Ç�Ů$�eݯ[��nH�%I��M�q�߽+������t�w��#�Hu$:�WRӶA��Հ��V�����=� ��|�7��Z�{�@bӅ������mߒ8ۍ( E}��?c�+z�pA������X�tX���K�w�/֝=�媰�-S���g�0^7ht���^q$tb���j������`?��*�ݯ���l���k��'|u�k�۪�����Y�MG����i_�awnPP��^ Nf3�֪���A�H�b5���'^p��B�;�>>ҽƾ�������&��Fl�΁6r ��q�6ހ��5�v�񊯢��tm5"]!-B��W�<�3d��:6Z2������=�*Y���#�@;p�����g�~��r�l��\��kUl����h	E�=H9�<khH;E6�&�R]م'�W�Gd���ݜ���
K���=h�c������B1�Q�<���[�XM�^J�>�S^F�b�랹4�;K�8�8��X�t���������|IZ��e�?���\�Gr��>&+_�����|��/��i�Wf�p��VwI��P��k6��a�$s��*X�������L�X�C��F���I�G�r�<���O{x�NVX����E&���k�+�|B&�6z�*��+���S3��i��`�?	FT'0���J-�1D��I	Z�����C��Mywo����@�I����@�ju�����ޙ�����r��HMt�����D��y�a$V^	�(��[w�ɬ��T+Kc���!�P��~�u��Ke!n��m٬>���N�Os�)�(��l"�}�H�#S�S�^�̤��ץ��D��<��ū�ؑ�&�zf&��O�ۈL���",�U���[���ں6����1gEB�5�"A8"�y��\' �G��/Z���0��Ȁ��ø���4$++�
u�$�6K; ���+�$>?*1v��@��	H���W��*��޺�,o$�%sܖg�ekQNqQ��8���yr���.�$sޣ;X��&�zm�3��լ�d�xVX5[��㝛�{ҎdS$�����N�xp�N&R�R'�l�Ɔ��[w)��b����i�s�=u]ln�lZ_I+L�B�"���g�:{~���=�o�/�~�%~��������u�AN"�Ǔ���g�"f�7\ ˶����V�4�����{��Ғm�h������A�>=Z�7S�����M_e�X_��S\�y���naH���Y�p�ͪ�"�o "���,�T�C� 裙CbҦ(/HԒE�^$�*++�"����nݺ�wGy"v�7E�7�Y0��=J��v�l� y�/�$N{A6���d�-�p��	þ�����'Y!Q4u�sy��Ƥ��;6�୰�=�3�t�]_��B6M��沰�~|f"k�����-�:�ࠒ:x�}f�V�t�Nv*�ͼ�R*Q����4Q�0q�+`�F�`������츼4ʳ+n7�?t<�,F����ٷWc� ީ�Y}�=ħ�#ЧY4�]BB��^w��Ld7�t�A�I�3'�{�1)����7 �Nlp�i��%p��55�Gڒ
E���M�
蚘��sW�H9�xc�Ki.~���2.L��ϤE��Uq��_�]�_��*9Ǻ�A7�{{�γ���)	�~�5w��O��_�QϦ#:�.�#2�X�Odڒ�װ��Q�n4�m.���e2.��z�\k2Q��Q�����1~OV^�FPg��Ʃ|��g�t�� b����}}�Rx�9����p�
E-
�\O�n�M��E������
i�Qjʓ�#�����4�&1�Ҹ���ҭ�x1�q|��+�'p��a�ϯ�7-i�������Ԍ�X̖N�t^����Fs�te�1ϝ��{�2���%Vevb���@�alw� �oW�i8�tܒ��^�&Cw��R~<%u+`��͒�+�\��z�6���g������;��K��;���[�.�2�[��&����;P�I#	Q�=V�2^���Z����F��y�>ܶ�fی�bT�/�nc���u�k%8K�ۚ�x�Ǫ�P���H)�^w���֜V� �aܥ���n��������O"ϼd�G�_G���au��{ �5lK�h��1��� mXW�~7�k�d*^�`�����.��'4V�:*ٕ	J+ܞhɖ��f������d�_� ���X���u�셣p۶1fG{Ф�A���z!-��E<�ʖJ��W�sɘ��߶�q��9����
�95��c��O��]ڏ��䁨��
��_����#���Ŏ��<���Z_�a���`G��Sx�p͠�������֏�A��d��8�{nK�����\4��:ʸ���v�9WJ[ ��:����C�苋
�y�!�P�~�
��nu�����Q�n�Y��?�����v���?Ў�QC�o�E
� ����ٔ]�o�VHRAbC�������(c��)�uу\/�״I4������
�S,�������>1&n��~�8.{84@jѶmUֺ���صI�����0�����1M��Q���Yh������#j#�BwmbE���T�CqTY���e�q��q|�J����&ꅫ���.�xɿ��K�M��!���Z�웭1k
��Wii!��2�����U��Gr�⧲����;���_���Y�WXm�~������ě�||෺��u5���_��Q]��`Ƶ���O�Z��y���}Kv�@�n))�Q��<%�xk�n�c�[ճ�Pwk�+ZK�~J7p|il-Q����ufT��B��N\�c�!:/�ͮj�x���ڂ��1�e���DW>C��Mu+�۰b�`��o'bN<��%���Fgը�7�[E�9Q��!�ɸM�p���jۛan�M�%��6��r]z�d|�^44jg����J���L
]�0?��;7�1o���[��Y�J��Y���LG��� 9�k�Pmwwr�d�K���$��un� �f�|Yv&&���?ˀz$ȁuh�����.��<H1c<��KI�IK���I!��	Q�����u1k�;��~�+�5p����e`I���p_c���h��6>�n@�.�͍H@��	?+.�m}�Ծv��� 1��r>��=������QϔeX܉e{2dw�N�o� �.�*�!����^��Պ�yvx�J�@X��/-�T:�S�	k�MҮ�fLjz�|)!�"JD���=��%��2L(���hYHR}+W�*�$�I� ���
�*i���	�l~A;+�?�;Bג㔶y͛�+Xm�'/��_����x�R��)�ޓ��:YM!�qs�y��[�-����H3�ro�چc��P�eK�geqHm-���z�)����YD-�e'Nr0
	�;X�Qǩ�#� P����'e�#n�k��{\��.b��E�5�s�΍N���+++�& +��X*U#_4�7�e��O�BђW��B��q�����~��q�~?q�|iM�D0����?j����n%�Quڐ�~${��E� ����2����e�ީ��uuJ�l�qi�z.E�^u��9�-���N,�!a=a?����ꅞ�<��*�vɋ���rQ��]��˥���E�DZ��������*�M���F*L����Ͽ���cr�r��m2�L����W�w��T�Y~�?��`~Y��s]AJ1�AOy�:�'Hm�֊:�K��ᖃN�������ql�,F��ժ!�l�W��ܡ�B���RE�iU�b�7&t�۾�=�6)���,�ϫj`v�6�~y�eS�p�����^�П�  ��`r������))e��A'`z���'�8�8�
a�´Oi>of�F)xrҳ����ؚ�"%�<@��{nlv�q�g9�pq��oŚ�w�1X�[��~[HJC�v`�0X�Q���>b��I��������q��, F5t7�M�To��Q�gAf�̽[��3~��e����K�Ӊz��L�[���t/j���bj��%&&vX�<AS%��T�����q�ױ��R����A��n_u,��UWȀvP�Cp�WW���Z���[�6,_��ٲ6Q�����(͑���F�����-��ALG�
�~S�:2��>Av������Qu��4;��w\�Wm7��I�.FY֚���o\¯'�3��i�f�m��>Mg��M�~�
�=�ة��:��/%��m4����o���?t�e�����>nlb�D�	}����7�XX�f�u�D��G���١�7��-�+lR��8�X�ۗ�%���������Q'��x�1�ֈ]��8GP��o	��3�y���6Ŗ���n���T�A�z%���?�C`����xUVk�旰�'��_ѡj��[�F:C��y��:ԓ�tA��[�pj2:5M
a����Q�EӮ�W�wom�G*��5���Ѻ+�Ќ]+ j���b.]'��j��e7ea�����S)�P3ʲ�A-Yn��K����v::V�Y*����):?�P�F	#��#��a?���h;�?�ݹ	]]����<��n�E����:�������2�a|������	(k���y�"����Ȱ��һ��h�9��Z��ݫ�X�4~�637Wx�3���y��� Nf>	���vz.��m�fҜo�Q�iɲ��V�b����/ދ	�!��B<I1�qo�>����gE�|�Y��O9�2��,��j�i��̝�?���p��QII�m���%��
+��,��U���$�.�!�tV�|�@Y�z�=�i�*�\ZA+9�8KYq����ݻ{صK�mh-b}�i�x�.h�b0.��]��X���>ͷ}���z���}�Y"�-2i�ں�ܡZt�^OD�O	��ĐL1��D�g�����#����G/Z�=��""�R��-5dL�k�-ݒ6�`��cz�PG�)���r��j��b!�DDEO�ʌ�=�P�<k�ʌ+���JI�Ũ��;���4�ݔ�ַve�!^����6c3���f9-V�ަ#�Ŕ7|T��,������ѥ~����fx�vh#x��n#����E>���m	b&���S�
��iW6=;s��1a��9˶�������f���0F|��0>9�� ����آ6Ҿ__k�dِ
+����e�g�E�s��dfmW��-L��)E��fx��q�&>P���<;�<�ag���E��Z,��5,��v$lS�s��w�C���y������"�Y��Z��)P#B)$!a)�oof�<2:G6<4d/N%��M�H��M����/������Dx��NOT %2����///r�x�:���i�Žh9�Z����i�t'g��9=�R�d�;PRZfP:ܚ��k�.�`����>L܌o�]$����ؼk��/7A�Ľ��zc�֙��&�����Y�[�9�RמvR�<M5��
M�쑡F^�_Q��=�j���x*��OM"�c�|��Mu�}�������XDMi�LYl��{4�[j���ё������f���M��=�?�R�$+(�hp��y����S�5�1>�3�q�~�,"���i��ؔ����A�&eԱBk��I��L\��w�����d�����e�嵼o;�D	(��@�( �Ć�)�K������Q	A�4WX�"�����e!��tpi"��v�mi�9������^cT��͙y�}g�o;:m�N��AǻE�����P]$(�}����̽�.�WH�$�^o"�\/{��5;�ݔ��1�ԃ}3�9A�_y������S���U�?�`W�X7��P*@L3���r�sK��|�w��eB1�,�exa|�B<����H�ʸ�v�\�2/XeG�a�]�������*E�����A�n�s���@N�69{�I����w�.2��c=^��~���ۦ*��НNO�I��|��J��Հ���j��7+����9ן/��Q&��!:2v�3�lVF�_�bP����'y]�&j�3r�����F�3f6��ʄ�ǘ��y&y|q$�jiBuY�Y2��7�r�-��7���^!�O��A�"޿CPE4N�|R�ը%[	�5� ��tċ�ŖD��h��`tV��~C��6Ӛ�&���\��6�։`��Jv�ҥt�=�MɵzdY3�@z���wjS/�����Z::�@4jjj^[��<1*�
"�$��y���ÁhI�� b�y�m�}��N�})K�����o�e��¥N� [���|��sd��цԅ.+���~���;|�4�2��"�}�g�W`�f�h!��؟��3uQ!(eW8��s�@s��̥LZ&ʺ�Sf�,���V�W�1�A�~���f쯛��&���.�ﮃ�Ի;e�ֵ>��聁���Ho���&���c�`���1��^.nG�������u�}gRD�v4�Ք���TB{�ޜ�i0fu�x���,vj�{_�ָ4�8�V��i4Ė�?ީ��Vs�����1hMf^~8Cr�f��	�����7�ѩU�M���]���Eep�q'�>N�HR�Ո��/����]����έ�$ˏ�~;���Xƽ��r�K��������n��|�������`���Ľ\��'�@��{��!��rUh5}�TGi�Q�"C��lrQ�cA����4f�7*4�Z��8!�o�k��8��^f�]�xB��jy��v�C��e�
���'��+vG�,�4������oG����40ٴ����8�/y����u�;��U�A�%�-s2��K�� �uX�:�������9]aN��%�0ӷ�e�[B���;n�K�)���66g��hͳ/���K|T�D4���ƨ>nR��6Q��wi~$��L}S�������`��Tw{{V�$�`y3���<��Yl2� �}X)B^���\�;,��D���_�[˯蚽��\����)JLkb6�d��'������c}�>T����JW�ʽY�ȹ(�8AX?jbi�	h�׋j���<�C��~;\�����y�>���A��JŲ�X�岍s��T� ��f���� ���M��?�� Ѵ!Wǥ�=���
W^,`"F77�i�e���w<e��y���|5��s���XT_����<�GHO�!�yq	��|� �p�<3�e�G�����eE,3	)��&}u�*HVZ`i����u��qek�$���p/֤#��A��49�p��f�.��Fy��ȋ�@4��	䢮��t4�[�T�h��y���/e���Sԗ��ew�/�ڀ���
��i/W��bw>�����+v`tR�ɻBg�o��?	�ߏʼ ��@>ٴ?wE
�l�+�Nj�BӐ�|�Rq���Z]�����ew�g�@K�7Pf:/��['wy��600�T�#�:d:!���v�+�U���r�Uĭ�S��oQ���r�p����AJ}09��?��7C�Zgq@6*��P\����[TD�8�e���E%J�~�UrNVa��.�yi9�;~>F4ժKQ�@��I����o�y�r�z5�i�c�?V��>CnsCfY����� �����J%��S���Ώ��!:A3��m�\G �Υ5u.N��z�Cp�I��9��@$�� ��ֵ����#g��)pm�$���N�{���-9p�$E�6ȅC��GK<{�Hs}��`�<7���ᬿ��x���ۏ��V�^�# षCn��;.���8�"��J�]$9��ƺ�k�:4es���)3���z:���v�s���!75�3�fž��Ͽ�]�3%c�箩�|�C�α�*n�\��9��~s�	�����/��V}�Z\:�UjuFEi�'�t6�d�c���ן����2��"���4l�7�� �����3�����L��zz/h����GSmD���X�������7��v�s4�I>���j�>hrӇ]@W��ի��r�ex‽�[��0b���%�|�o��a��� �cQ�,-�)?캩O0@�/�)�T�2b� �(I���?�����#x�Cp;t�xo��� l��Nq���2o!��Y�׭]�Ŧ���s�7#]?sq�^0�{t^7DD���"�����b�0I�;R��-a�+�����k^��Y�R���o��U��Q�UI��H�����;�vt������Ӂ5�J�%[�d6;��Fg��������)ڨiK*�1Ÿ�Ξ���;�˲�ng^t¾�!P'� E;��89!m�m�ߢ����Վ�
s��Yȴ�iND�I$�rL��P>5�6o@��|m�7=�?�m�Ww
�(-�����ڊ��9::�Cț���č�>�cH�4zp�x��J��,���2^_`fb� ޝ�}f���"�&����+���wG����ܟ~#db
!���eb�^C%�w6cA�i���q��2O�`U�QV_��/� m>r���@��O�.NQ�'��;;�EO$n���2�oȈNFc��LHȆ��zg��E �	I����%|mڴ��>I�+�Rp��1U�d`��,aԗ�z�t�b�Ѵ�-u����p}�j���͗-��7Ȼc�jS��	�#��&fSS��F��?L/� �Æ~���OZ]JF���.0h���<n�	�8����,���rP�%z������ղ)�	�y݌3��e�KT�v8�٩y{{�v���jg�igD�$6J?�=1I���m/Ax�6�z�֦�֧n�i�͗����3F_5g�.�S
��([4�E������ٷ�G1�	.o���G�;i� \�s��6�^,�b$�s�b)详:�O��n��AS'��ǟ��}��,���$+�e�;���L���@2�������Y���f�-.2FF�FD�
+���y?P ?�bw���4V?�
{���������[�h\Uw���@=�����ݺJ�r�5�ࣽ�u�=�/|jp��X��Ƿ��&*c)}ׂN�K�N�Y�N5ċl8j�d�����.f~�k#�nj��H�kE�D�*�=9 :����T�j݃R�x�����2�\E�D�=��=�gSuM�^��6<������]awz.O6;H7�6��� ���L�3�2ܹ�8>bv�ڀ��{�\z��on��A֜�q}D���8��vEZB ��݉�j�:��k���m��h	���N)Mz3��V�F(�ߦM[����HϋOH ��v_UA�[�~�(���-a��b�(Yb9+L�Y���|myu^��$�ԃ��G���{���;0t�K7�ۡ�ȮD`p~�����#���w��{��O���6������Y���g:���G[�����o�]K֫t��p�=�,r��w� � 1"Vj�0�<P�X��=ʹ�4wǡ���DVE�¹T{4�(8�ldjeEE�N�@V�c�e��NLL����6'}��6C-&/���%�/��U�7"����H�WV�чz�L�4�wyǾ�i�|�E6�Mw;H���i�;��O|���y��"�v'g���0��lmm�=z����5X� ���XwN��ӭN�!10z��R[s�5�r,��/���n�=M��I)�������rH�}}��ʹ$GlJ4��⢤P �����i���G����ӄ�.6��D�9Ũ��j*]�.-�@3f�hPLe��nX�Y��E�k�U������~��)*�)���6g�.�r �%�X�O�c�Ғ�*��ы�U٨�K��?Wǧ��YTnrջM���bۢ�L�
_>�A^{\�r������ݶ8���| ��x�{4kn�/pa��$�$��kp�ty�5��u�V�!nbQd;j)n��0`���B�o�o��x��E:�ɋ�ia�:YY�ͨէ�L��Ͻ�,Y��~�O{�9Y���ٴ� �{��? �b�������N�b*WG�jק���厖9x��q���uh�vjr@qi���o__V,I�l#:�ZX���_�.��5��A5V�zP��@��`=��t�#���n?�<��=� �_u{̆,�%^̡Z��~�o#�N�E�ק���
���H�g��������*�J"����4ŚnwoF{˳nO~q�S`C���ó��м~���{�؛����3v��v��[��w6��{ZG�>T�M<���Aq���I�ӛq�3��Dl&uH$NC#M�@-�&�VWE���;����;Ù�ن����<�9��Cgj�cPP�P|�����x�'��q�a/'���g�S���e�k�S�n�KQ��5��k���&*J�;N4e�2Ӄ%p�m��so7�pp���.fy�:����٢3hޕVh����*\�]H'�#S���ư���'����y�*���sf�w�"O��Q	Հwu>�z�:XJ��0���M���3�M*b���(r��i� �F�_�e�do������\�����Jpش�Ej0������B���rKu">	�)8��^��dfS�}s��u���uj��9����iv���%w�ٛc��q�{�%bE��{6>0?��T�m$��Q��)Q܅�B��6�����2�^c�5�>��I ��\��T�W ����e��Ø�QC ��͐(�f+T��B;w�!�g_��v���!7<�qM�+\���.Џ����'���9y�,Z�ӿf�1�;Y�oa1��e$��A��l�|=!���@2%qI����x���������Sh��p�F��\�T�x�4��&��?�9li2Cu`~�4����� �?�H�������
�K8���x��7��w6V\9nyEE�\�G'O��hm�� �-	׳�rGЕ�{"q�s󛆦r�������#�?���=����oͷ?�Ntiƀ�A� �b��?;��dq����-rqCܺ�f�cB8�'YC9C��v�An��!C##~[έNg�	6n��ľ�8[W��������#�K�dhK;M7�b�Y�Y�Ƣv҅eմJ�Ċ7����ϟ�� ����cW�!#5z]��>�8l �0�rX���A�Y�������iV�rrr�|x�A;Ó�I�e����>�Ian��ISA|[wu�����W��:��\tQ�w{��,s��Epu,�)�����Ę(�_��+�g��UM��Il�M������6���q��ѻ�Fcy8�o_�ސ��@� ���G�L��[�z&w���~ꁲ�g�N���2��HѦ���wxF�m���5�qxI;o��ww��}iqXhVE�`f��\*<JK;D#y��gMT��FDlω��� Q^1��@��%��|�O-��f���S(,G6���h,lO\ΟVj�86ê��H��+��~{='Y{>�����OO����f7�)�]�+F���,��w���B�I������O��I�urQ��-�IY�
�Ժ�j�|��bq��@��l�:G����I�ے��� �o�d��(��ޝ���)�Q(J����a{��f�+fK�C �	���g�֮���Oۂgր�^S��7]�a�<Jl)4�5������y�����A�:)*�mm����=-�������Đ��=S�~����a���hv���l�������� ���U�7_x��-7�,�fҷo�W�hf�-���7콧�~�DG�s�z�QZ����H{���!��"C,)��=��ٙL�����3�4f���^xt}V�8�g�n||<���o�\�*N���l��9�}����q)}ˊ�Y ���u�do�)�q`�{칭j�e7�������5'���\9����VhUT� +�R���"�+�%98��N�C��15�$tpR�>�:�ﷆ����T]����r����^�N�D8�����ؕ�{�&F��h9�����,�?���d���?�;1�{W��������p��	�V#u�pw����սϞk���Z濼83���Fz��{�"��i���+H`S33Ņ�d��Ҁ�����4f�f����`��>���U} �zuK��fW���:R:�.� �k*�Ī��?��h��[����-�B�+c���MJ�+�`��C95��0�w�N�	�KQQ1��y� X8���|4�
�m��Nokiy)�Ç�V7���$������K5lu�0t �OVQSs'ے�t�hB��ʱ���y;�N�)��oP%~���?f��N#\Q � �y"~��aY/����2��(�:F M�ۨ��������"=�?A�
��Bh�	�����:��@V�v��@U�(��3��������OasL��ak6�yT��)\�Xm-6��E�U�x? X�-e�/l�A�K��.Z+H)�
�p�:��V������"!��K_@�$�8:;_BK��~�T��~A,��	$�<��D�>�A3�3D{*�o���G0��z��-���n`��|6�P���_�!24I]�8"I��3�:$��4�}�^@!�������^�~�W��ֈKCx;Ͳ�1L d��%s��=�_w�^��� ҬT�@9���@�xw�y"�����	��۹��d[�N]tR�X%�2�m���F:��b��(�V�)�9� X�NS!�N�v�AU�c�����VC�)n�7#<䞖��-;�&���#s�X����c@�8���?����zu��#���@H;�#Yu�`����&�n ����2ȼ�*7����o?�z�ɾ#���,��_�!�V��8�F
X�'h~=�J~W"o�L�㛇���������������h�楥�TjD�[N�䎎�˸@OO]�i��V(���1D��>ʹ�z��B|��n�n�Xw�������A�s+�,�U�W��L:,�i��n2�l���,8��\��} '##;���]E^���)$�d+�t%��¾�̵a����###:î�l���4�\�������]c@� ���T����~}�Z�q|
DVOpB��HC����lp5�צe��*q�8
�ë16��e��-��Q��|�m�)��M�5������&wc5O�rJ(]H�F<h֊.3L"�[��zG睉��tO���t��|{e~�#�iYW(8m�r��d��2|��1�փ��o�E�^��_�56�l����Έ`we��?\9��1%��X�
q� DnAW�TMG�x(�1��|����D"R�J����?���r|�d�d�������tAii0��S�M�Z�3������VT�<)��I�b]E���F�����p�;X�@��`�z����:D���~�`����5�t��R����� S�έ�R���Q�K���U����	�T�I�h8'8��_���؂��I��-x�@V/' 2
�z��R�>�b0�OZ]�}��1S����t���@*0D����3���3xy�:�*h��j��"O�P+�^z��&^~X�>�����d�-7�W���a⏫;0_"Z�<�0�&w�!~��N
��ח�p# �R�����񠆮Wrm�^���˷j�r�d�����L� ����3��l$52��*�|�E�r�����C����F�"�:���zz��+��<0�
�u��/-x�	w��Wx�+��O޽ws}VS�O�O�dq���f��bf��X�O'���D�lr:����w�1�t}�%ŉ�:�M��/=B�h)iK'?�W
�E0�;s
~�/�fߨ�$n�������#��%�����K7��.�P\���&�/�O��2Y{T�l�����ky����IM����}<<~:�Ϛ�{4�6(��R�6�4��Y[��M��~/]l/ŷ�"h]_ �r��CS	U#�^&�N���Z�?��cvD�s+��5`|�Wr˖S���/��q�V�ˈ�Y��#���Ԥ��?�.�nz���������S��b��y�&�ɭ[���,�_J�:���jN&�ND�]�K����(������(RYʺu�CYk���:��^������\�:�0q���yȗ��z)H�{���q���03�&�3ZʺG/tQ�<�.ښ�VK�'z�#��j��~�:�R�0g�x�y:�2��H���V�񞙙��g���I�d�A�Q�߯>펿+�3ZN�9w�6���x��ف�G����W�3��[� o����)�E�u��4'c��� �f�S�z��:�_lMX�e;#膙� zHA����78L��-b�LE�:�d�h"?������I�%����ơ��ټ�	�z��3lںm���OHm&��U�b�)��i�Z�m�ѯkyG�N���m{T��&)���5����D=�b��_��Db��Sʫ�gA=�G�v��ھn��WS@�7x��9�!��j\d�����P^*o.���'�w4�=7���Nr�_3�k-��"׶-`Ԩ.�-��є?x"Qxg���A�6���J
�w��5r��S��ju�=B:����Dr���%a�;t�I��\c��{���Vڬ��ۨ�KڎՒ�[�Y��N���������叔w�&�+�ɻ��4����H2W-�ic����H]x?5D�n�����E�K��9�,@��^\\��ٚwQ��	�l������S_��|�n���o	��~��2�>�f�'�����+S1T�a�p�O��j��M{�*��g�b���k����4nu�WL��HE�pi��`�H;a �'ߐd��a2b��/��@ ���39��Hl�OBůP�mk[�ǭ(���3���e6{��gnb`��H��N~�+��@r��$�3s'��l*��$;����W{!F%�oN�����m�U�s�HJ��@l�[�8����6߬~\z=љ�3=lb��MJZt��RQN�"b{#�P�re���;Z�p�J� ��N�8	ڴ�I�$�?ӛ+�V��J+{�T0ʙ>U���klQҲ�QW`�:��c�H��X�o1�s�z:x���+��|b�ٚ�|�Ko(�2r��m'��O27����ǢB\�`л�Н�_�_�ё��U���d6��s�5���I))��k���q��M��azd����5�]�5��f���^hp0��<]ѢK0��Hc-ͳ���E��ˆ�A��]]\����su)l��t^��;�R�3�`�驃du���;s]������7^�#�Th�f��=ѐ�
��d4�Լ�a����aJݿ/?��\�:�S�{hđ�?���}'�n�D��-V���ke�E��i�\�r��?>Y�MO<!�ZnH�B��������ʯ���%����������h�]�[!�L�x.8<2�[���;�g��#i��Oî�"5��?�NX�%Yr{�|��ASiB�q��V�MU�^�0�-(1OMME۵��>O��bA�m�{�G�����սyG�i��#���.़Mޙ�#�p�ĝ�â�	G����'?��废�f)lF��d��M&x��f���=6}��sb0�@�ܠ�K��ȟ1jߢ�(���T���I��M}BS�Do� ��>	�w\���=�B��m��w��ȘWnZC��3��oy̏ޭ|t%�ޘ9�h- �@�F}re�7'z:&��3E�`�o�w �Xj�Yٸ0[c]�#�Fr�*\xy��?V�c���P%�-���04�"qr�mn$���Y�>�w�g;u�b ���4���B��}�~�Q���J�v|_@�Fp`C*����:��#����|��n��8�3iwM���#t� �Nȡ�ܢkRƨ�����k�sO�н�h�j�����vo�.g��N7����}�}�.D��B�|��/s!�W9��- ����ۢ��g �����^ ���z�dhh�3ѧed���7�PO4h�E���\1��L�b�,C2ρN�}{F7g�;�ߙH��a+�:6�B����~M�uR��F���L���)f,Y�n�e��FQ��Z^+��P���5����̖J����'���7Xc�-�j�d#>sGU�B<!��AK����hG�,�o���cEm�,�D"�'�v_A�=�n�<;�F���$���|sU�v����'��J]}�ؗH��Ķ� ��Ĕk�Qvu�G
�<s3����2�L�s+�8iz�uk���T�`���ѻH���vn�1X�> f���8�D�}m7<�&~P��xª�^����Qc/
?����д��=��>W���4ԝ���3����z������]�F.\Ȯs�I���`r�)=���դ��E�y�SM��A*L�E�kĢ�����Ӧ������\߿~����X�D��C3�b�H��䃨r2�hϮ_����n���KT���0(�JG�F9���@���P�ɼ�*|�8��X#Sti��x�zC;�';>1�ۦ(����[��Ϩ�}v�&�c��_�$�D�UX'R\��o�G?�=���U�Qk�آ�.���y�Ψ�	}2zQu�yi\/kj�����1C���	G3�F��ݡ���P}"�~�
�n��G"ɯ�Onn|��e�!�F�����$dJXb�~��s�t�K�w���!�[k/�QTN��e�N��Ie<t�Ӭ�[YD@���:����8r
�s�gx�y
1?_j�:�M����,��^�h��?�:2����0�GM̚&�wJ@6AS�!Q�֤��ۄ�oõ�o�����V�b&��� }8��3�4�������e���z�yM�KS&_ְ9��5���f�}έ���+���L���\��y���HM�{ZU�wKo��I�n������h0(ɪ�ن�'�_���8^)�5��)��5�k���������
H�'Q��M&1�ք�E�{N�5E�ʕ~/;�1��ŶY%_ N�%�81B8�z�Ç:I�Dz/)F�����=P+�a|<8?%����ϿJ�zo$aǞ��G�~(�FusO��}�"�����Mr����lXɢz�^o<��8D�(*��O��҃)��n1����t)�������\՘<EL�Z�����d���y�eHsͶq�#�#�||��'���Tv���T����U�竎on��`0��F��S6�.{O�n!���;U�T?Ő�
GFF2[]x�km$;:Q�?���F�j�q��޼�l�n=txp�^:ڞ"b�n��q��6��[��2��x� z�G�c>Ӟ�� ?d	]���H+�R?|��T]'�T�N�v�Xs��h��S��)Gx�u�m��u��E��d5;I�'�U���k d��i�#�S��v􍳗��W����,���TL��W�YQ�8g�=�n!^J�����`���b�%¯��)�����:� ���? �~�S(��y~��(���wDL���m�{�$d��<,��3g����V>ו������.�_����~AR0�={s�G��J$;13+P�$#���8�]�_�1�Kڒ8�����z6���˪�dk�	�����wmA�iM._�F������.(&������|Q��ebbb�[J��}t;��m�ڴ�Y0���@|�mҹڕ��g`��3� ˻���5�Y�YYb����42����ZH�R��Q'��L����Ǐ?�L�q�������曈'Ç��z���UZ�.pF�u�Pu}��n?L}ŕlǓ+n>\w��frc�&�&�v'��(W I�p�N�3#����ٙ$��_v#_ܲ�q{�{��%�������/�,�؀d.�̻#􄬬��It�����d����m�v�\ݕ�27E����:�e��ݷڐY�Ҏ��x�:�0Ā4���IhJ��W��W���j�E�������`�S�����W!j�Q�/^<�����ص�߮��׽�=�j�
��������<�MB/昞6�L���YC�H��߂Pp��o���HF%:J6����G���
���-\D��?����$v�Gǧ�ݚ2�ů�ԩ����ฏ�y���v�X�n�߸���ZOMLLlJ�&�������恰�8����.x��r�?n����'��nFS�_UWe�m)��z�E��jE���.�gzI��D�o�j.�?�Ou�UV�X �0j�ĝ�J�1K�Zc;f�{�H��7�[7�Tla'�����
�ݫ�r�>@����Q��(_&��q
Y �Y������b�:�{���� '����Mٮ�%���Az�m��M�"1�i�n�N��STe����'3�Y��
������l�$�9�=C5�m���^g�x�#��<���?ۀ������b�7�]�Kv���f9�¿G�#Ď�-���K�ޭ�4����6�|7Ch��Vag�<�RY�r*8H��_7��>�G��H�C�D�؂K��K�O�9o�wD�a���/�B�[L��R)�T]��F6��h��c�B5����]i39GO9��+��hW�̎��9ŒӤ��vH��)�;32��mS�3��U�����:�:���ڵY������)��l^a� K2�rindLx ��2.��A\[C$��G�2t2�����2�}�L�	�����#� �UR�;<+{��P��m$��GBΆ�'r������_��&�g(')�cD4�����V�K�R/��w�y#Vj����56�G	d{��3� ɂ���Ӥ�*��tDs8ƓAsE�V���Z�+�t;&﷘��|c��gQ�u�U?�5c6(���ƋP�����F�翺H�35��B�M����6���o���;+ ��nf|���4'�`U�=>��yO����I�^������ooU\nB��U�SJ��l��!�I�(�f{>f@�ܹ01 �����\��Rv���%mZ�]-���)���Q��ؾ��[uuQ�>y�~P T�4P��� �C�A�}���a�TPX#�a��t�u�Z��q8��rl/Sݛ�E�h�G^PI�m�=��}�u��|��O�t��ʓ�>�=������c�.@LD��y�g�+	���(Զ��vvvwTT��lXȽd�n8��~��z���� A��+hwEsr��"i����Hw]M���+QmvAxMb��V�dj�$�Z�me��ܸ�{�}Ɍ^ B��i`�1�W�m��)�+'G3�*��fJ���B��1P(��r@@;1�/��*�>�� g}��d'3���q������/�)v����@��СN33SSS���ї��4;�/��
M���}mm��D�j��Ir�D�F[W׌ʹ��	?P�Fy�w+e���jC�����"���78����z���7�Gqh�FN���*mb5�\�q�����0-��)L�Y�ݴF� ~3Wk�r#�F T-���l�w���X�M�ᩯ"wo�Q�;��T�s�!����VX~�|:��z/�c��e��֢���:eu����!�F�i*�O^�<SyG�>����=�I���cR� ���}�iփz�S+�������k��p�L���N��
���m�E��=���U�Ϸf�#�'\3a�����1�(>y��*@A��b�{[୦:ikr���@��V�'Ƣ��-9�E�nC�rY���tq~�iU�_�*�̩�)��4��ֽ�s����4���Ǭ�7���ۯ��.a�L��D�޿�;�5.�5hgӾ}��N#��w���G���@3�Ar�P�����W(~^.�e�a`�wI����C���KI���tc^�
)�ي}/{��_�u�v�'A��t\[(N�t~�M;����精nD��QPJ��τ� �J ���0�ۡ��4кwuO�=V�-0qKxT[�E4ө��!�
X)�Q����_[qu�~w�C�Vȅ�3��?��J0'cQ��&���ϻ�N�M3;�{�t���0����%J~��cu	��c��t��r����v7���C�BqWX���+=��߽��*PDe�!Z鄦�E�#Ĩx��i��R(����t~5@S�)CQ�!m��쬽=�^�d%��
�'.�(z,��(UD0�ttw�'.��	GGE�}�5�(��٧��q����ǤP6|m�r�K/0h���0g���!-�w�}�r�ˇnD�������(o����yM��!�}��,<v��R�c����DT�M��q
�[�(���m�q����3qmd�M堅�g�G�EӁ�N�?]�l����������iC�EvX,��ڸa����(w-ӫo����Kc��X�_�:�,����<"K�3�g�U�Ǯ�[]۠�\�� aA�;J
3n��&'��>@�5��% ���(ɏ���}Tٶ�]��d~^�X<����#��(B�)�.�>�=�G��j��M���� �55	3aN=�FH@�5��%OقGਜ਼v
�~�o��>��}�0�wp�3&*Y��o����{">����+�o#�L��GA6N�Ȯ�=x*�@l�(q�.;+b�'���:3���D@ ��F5�t��w[utt:HO.�M�*�r��l�P�,�{6����k}t��(��.l���f[�r<�/��j��Fz�6��������5�U�7ڝ�V'���55�A5Q�F@G4��>���a� ����o�:f)�����H��0�9e�]P�e�-��:Z����m�we�Rl�9�[k����I��0�훳����<�C1��hjh+�'�O��P�)!�	��j����zߥ���CJQ13��U��a�Kn~~����qs�,Cb~~�i�� ux�銷\�CD"p��|v�$��XS�6�7Rz���(��Q��Q�*��j�P���T��z'��@�(F���0�a�������H�J��O�g�˄����'X{���::|�a.�_-�)ֺ�&��Rx�PZ��� jr���ݯ+(˒���i����i��[�9�mSr���I��ұ�ܳ�rI��_ Q�y�iٲ���>�%I�̧�g��䄄�DO7Gpo⛹��Ӝ����1�r���������/���^�[����<��a)��9Q����L��穝oШh�Zq���<�U8L�]y�<d����Jy�b+Τ�T�ڿA2�փ|�k,-�i��j��⻚��\U�����3S��Y6�Zi�����Z���3L���Ԕ�i�{�; |�����\<��4Hg ��+�����"l�
�?s�?V:4m�*'z�h���O���M�e��<��y�"B�t���{p ΰ3jU�<�S\�j̘�]�'��c��(���<$h�}B>J00�nY�]�����+��smB:^���4z_�,��<������G�<F}ԩ�;H?q��O�l�p��#�Ϗ�RC8������+��`�JY�gJO����3hаl��Ï�;�d>�(|5p��T��Օ�Z��c���Y��Q8��#񢪜���c��p�����1�TI�wd��h1NO ˑ̵р���^���L���P���0K�k��jf�3w�®i�	a`�4�
��vHS~�.2�"��*h��|m��
A�-��m����[���ޥ�"�1�
.^/ ��S�m��D-�i���Uc�hl��z�+�VO��{p��rn�~{���3���Xqsz?Hy��X�&�Y99:���̑�Lsqr��I<�y5��V߷�0:*S$	ȡ��4�6�4+�J�c妊94�6y�(W��`.-�����'u�]��g�:E?>G�?��1�v�ڐ5~�.u5O$j�D}B�tq1��^T\�'�Ј-*榥��}f��ťu�]�G��.�ʼ���(/3UD��_"�F�d�t�h�9�����Ox߫P9IF�����B!p����N���5Q��̔�J-�@u{��H����Z��p���K�P#�)��
�S��Ǫ�=mx�̴�(A2�CV���F�`��[��{|t^�!#U��	��`��)�����:cc�JX_�ҏ��U����� �⏨�kVڼ��;]O�����d��N�[�Kud�p[��y4�$qwJ�/���������E..E�;r�ƞ?(��8��a�ը� G�+mSq���X���y�,ɑ�ϽHI�Y^Ƕ|~vq�l��K-X��H:�E����P�����j��TB���b׵�3���NLLl%Ek>yL�t̶e�+V�UX�B>��+�7��P�.�ܰ����_�a���R�F��(rϛ^L��{�?@;�X��El7�� ��j6ߑ3����, �t�d >'�*i�K�Xr�O��QUu[eqR��x�����.�q�8�x.n���Θ�g.4���ޅ.�J�I�m�}w��BQtnη�LM�������9�m�b���@Uf3��:H���W���Ɍ&�HI&xAN����QG��TX��g���:���St&'2ʯ�������k��F��_��0!*�Y�ޙ�O�_Ir`؋
��ziz�-Ŗ�^&�G��o[ȅ�K�,]^
0�O�<l}-^��cE�4nUĚ�_]绡Yf�?�BN/��#^�������b*IH\G����[��*�O�7�a������窋 6T��]�(�����f���+��u�
3z؍t@8��V�����ƫ%��{-�W������~f?*V��?���h�x�#�����nT��7�LAA�畀ھ0ci�l��#���t1׳e��=�VS���y��\�gQ��-��vd��7SZ@�h�����O�VD�����B��!�8�ܦ�2�Rn3�3���gb����S��.2S��:直�栋�@�Sϭر�w+	(]��� �9A�MDQ���.#+�3%[����!+3���%TSӛ�&Ac�������N�{����ﺅ��~��؝����uu
*���Y�^����#gQK�pr����b����k�:Hޖ��=�?����O� ���!g�uv��y��y����Lt|��#:;�y8�ޅ������@���HT硁S��F�b�R��� '���4������鮨�gSuQ���_�v�NY�,���h)���`���!L 8]W�p N��
��Z
����+�(��;́���ɬ��P�N/�?bv�����Q�(�<��s�<�T�9�%0���)�H���q8܁�E9L�l�d�K���d���|���/�!�`ݬ^�`���_�����RԊ��ݜ��_�"�[#;՛#��xY�$�>��2�ߺ�����=l���:�$��f�9�P}���Pٹ��N#�TG;T]9��7�m��_����jkj�ѕ�C�F+��i�V�e�Lg����K�BAN��fH. ׼��r�H,s�43����;u���j�FF[[��R�U%v����#4�����a��m��a��9��񽽶�s�	����t�49Q�%�}��AU�f��
�UC�|������� _ 3��Ё��D�U��;��p�&t� eYs�F�IP��Y��f�,�T��� <�C�D�?����g��PC��Z�&�ۑ�˅��3st����E������=K�]�Q���_��5�˗O���#���I��^tt��ss��C�D*�ڢ �)�c��sQm<�l�fb��M��?n.t�@�2Ƣ�����spp�V�V1{�7�T�5���oF�����T^l�
�H�Ҝ�^+��a~*G�̧�1�|%͑-��V00��y����� �L���_�m�}�T�u��|�2���ւu�����<�
0��&9޺ё=����?��E�!��c��rE��6���Rr���[��k��̞�KP�1�-NF1�G�]�#���Z�"�_���9�>\����>�u��f�Z*���Wx!�]���έ!�4��&ŕ�2x��j(���~��*�m^?�POQ�
c��^�v�Fs��:�שO�H� ���L�n�n�+M޳�d��/�s�?g\t|���?�P�XW=<�̈�7��eAB�� ̙j-/+?��߷��R0����bcm ��ZnF��˪�����>"�
���=�;�Jy-��ˆ�����j�\F0u'�1��=J�2�c13���9ͯ���w-2�I�pn	���
t9t�[:�/;������1(��-�$\(˳�rm��a5㮏�������}��Egg���[�IH�'������+��E�G��$��X]�HJ/B�JJRC�4����|�-r:�)B-չrqX^k�2/W�|0�1ŀ`�R)�8����mA��^]�(�P�HPƅ�V��_��#�H}�j[���Lt1C
B��Ky�S@om�71m�4%�.�{��j:f�gt��n�dK��D1�O9�j%�d�_<1��F��Of��7���ە��@�[�V|��~�d��c��}n��+��c�V��:�á][���|b�	�&}>�쓠a�ռ0&��e��^Y��3�(���܃&x�ʹY=��rӪ����]� �@pUƖZ;���vЅϣ$��Y�����;>>^ZVVv��Q0��5�`_�EF��M��>.��ZtM����'��[I����xD2zz�7|�U����*�Q��z��V�q���1�r�`��ϯ��R��}߾C�~��bN�*Ķ-NU��3������.l���3*�o���(7��d��I���9���Q�k{�7o21�n�xb r�vF/���m�EEr�����Ӗ���*�Oe�t��::�i�u����n���-��}:H���ڢ�8�;�q>�4:<ꉰ��������1TV�99Ơ�f�0c�_�oh���������}��Mݿ������^�u_wC��@qǬ�#������*0`���_"�1Wׁ��f��V����:"�����Xm,�$M�p���|/��N��;�I<���G?`\��3R(�^s�*Cp��q6¤��^Dk4
�(��[�ga�ۋ��Xɞ��{��,���i-E����D��#�u�:��쮹���d�&��Q�����O��JŽ	� �C333��B�MOORM����J��ڻ6���[�"k��^$)L鞯�����_���c���#�q�l,�*��l�-1���q�Ґ��!4fN,h��������(��Z,Ƚ��!;񒼌r���XdR���m(�8�uyΜ��tͿ\�/ЯQy����T�~<a���v]����'䴵��.�V�}��zl��� :幰p���������phcC�3C���a��AY�:������g�x{{m�6�ı�ǡ�E��OzF��꛷�I�L"��;��1��7OT�Ͳ�_���,��J�'qf(0��d����j�8�1��|M����葸1�X��6��:������(��N��ِM��.<�����ۈ�h���a1�4��u�̨�Z��2/��a+�Q1�BGeڼ�@%D��8��>��i2x|Y��o�\�����o���g���@��趒��gz\g� ;Q�o���$�D������7�&��s���9��t5��F�m����U�HK�
�v����[JC{P�M�L	ʪ�^o�D �
��d�H�ظ�W�=u?�Qo�`��_Ww�d��U��W��K2KC��)��=t�yK_J�W�G���"T��ϾO�~�M^?�<2�0���X�3��������gY���,C��0g?�[��H���H�@e-Wq(�A��*X0�+`��� ��`��m�[SS��� ���g��^�/�36�m�@<�/�	�d��l<�K5�X��S�OE}qz�sǋg�2׆�:�%���� �.C��]y����=�ﵪ�]�+wAJ�}��?>le�s�x]�݃��O���憰�$�^�u��#��:��(M�}�F���mm�<o��5����-���ţ�L���Ƕ�D�+�F����k��S��Xxv���Bbcc�m�u�-Qn�@�V����������=D�}D���k�;��	 ��c���w{�xax����y����U��@��r��J�������1�Q����9�%���S�o�i���v�� �6��M��ktMD�j^a���J
T�e�e_HkpQ�_�L�n,K> �^9�/���Ұ��f�W��Smr���Ԭ��/��&0�kH��kj��NT����k�QŢhz�2k�>�G��i�&lN��65t6E���2�;o��Y�p�\�D)�wٹϫ��#!��R�G�N�Ɍ�v���ut����K	��zf���Yv{}�^wcZ��XB��1:�!N��jq2%���]���W�Ex�>@�٭�J����؟�AW���?�����,�>�����gg�v��g4�۽1۹K:�{ ��t#�~�ob���ǥ/�Ĕ��]�-�]b��?�
X�,8������-����@�	����py���c���zu5�kh4���wW���u���N���x}���Z�L&�.D��Y�+���r��������-�hx��E.nbkt؂��x�L��z=v<5Y�.L}��E�6�l��f�.��p�P�	�I�Ϩ����g�o�/��Ӷ�ң�j=[�gS��೙��Y�	P�Mwz����g���ݯϤH��T���x���p<��������˔�Y�涨0ԂЎ��2Q�9G�;U�}Ʒ�<�09(_w�'�=��n
��T2�P���bt����g�i,S�Xc�����jD���ȦiI���W<���c�P��#?H������G�����;q�3�t|@@�G���&����D��]?))��$�X%��o��X&W���p|���&0 G�OWQS޼,c+çk��ʬdS�X/*���%�{�`oxJNA^���M�3;�WO\C#�es������N���~���qw�
{�����y�nݺ7�(���t�)7�E [�P� �w�Ve�5X���m�[o ��5��US����,�L�;2Yx��|�N���V������N@ٵy)FKo�L�8Z��O�N�fA�����
��?ߪ~�!|Hmr�v�yP�掎�yZ�h�羍�YU'R�CKϞ��Rn�^�A�9��xJ�9k��/X�FM&����J��R�[ڶ���������W*��4�Z���Yʶ�I����{'�^XHw��(���,��?��ڡs�e�i}Qu�ڑN��������hs�-�H�h8�k׾c���Z�'�����19¹��V�/�)�b��[ټ "�(ƛR�wu�M������{�~� Dܪ�*�8�TC�[ӵ�}h�.�,!MߗJ�ɤΥ� w_�Q.����?��Eit����,M�C�3��g}�&��G߯ڪ� � e���yP�m�������W����v�W���~��_[�.LjY5���`.����gi}������-uuF�$�5&''�F8&�kM�@6����lmEw*5�?�L�4����u��II;��t �9���� |ۆ�� ���Ȼ����*�!��T�X�+�� �
���p��.�V�^��E$�-N��W"$���V���.�9s�������r@BK[���U+�Μ.R۵kj�̰-�ɶ��WSK+�ӊ��;�3;fgƱ�Ɏ9���>�≐Ï~aw-Ojq���8����`�!���4P��X��^W�U~߇���aM6�w"lj��W
"�����t!P���\�>�	>�����ӧ82jdFi�O�����N��\�� �H7P��\�?�1P�;�4�^*����9��̌��hd�7� �Ӷ�O8+����U�X�gA�+q6�L+���T�֞x׬���8A�BQ�s�~�bkw�Z���P�ێ���MjOw�5�����Ig��:�2��E YI��C�@�6z��7"�c��� ��*!48s�Opbt��/M�|��r(E=66J��ݗ-����-]clmi�r��ϟͺ�n��̧XOq_ ��S,��=��nܸ�eU��E	��/ ��i��D��Qͭ�"���*��4Ν ��I���q�<
��77/�;0�Yuu�m���l��.�Wڑ[ŅjoJ�����43T+�H[���Ç�t���[�퍩�~����� ����*�7���q�r�Y�UcW���%�zPJ��>���Z����_��NJ�,R��-�����n�\)6դ�gd��S�[��BO>���"On�ڬ�#����������;G{y�q�R�����B`Y�Ԡ�f���O	�-�k=k&����~6-_����\�P���Ww����d����O9 Zl�
� A����n��_����� ����;�]_�6̤��o�T�1����cGX�����Ű��y��/��%�{(�����Ft�Q�l�՗��e����r.d,�mt? � ���Nnq�������c�"�|e+@�#��9յjM��pV��DW$j���!.���999��o�A�����hT���s����nt	����qa�Ϳ4w�:�m.��I�+��I�`ٲe�6�h��F<ph�8ݙK4�	��Q�)�Ƶ$MFOO2���;}�H�t�J�!W:G��s�Of*���}��kvFp�~ױ�l��I�Y��ǹ��E�7JQB�����dv9�����lRO|.�֧+�۪�!$:�CWN�^�G��|�*o���I<�����>�#>55UxJ�٬�^9P��}?续�jk�&���j>'FE��F��|�ɞ�y��8�`�e^�3�����nf�#�8T^~�[6E�����;a�6O���q��{zzn�5j���dV&}�DFT��NU�����8��O	rD}z����b�H�ڒ9��\=�X�-�������Y��W�����1٧���e��!|�w��UG��6!�_�n�}
�s�/�Q�;�~�@A���ˍܻ��=xt�:��(���;H�g�,�d��lq*6�(d���&HҨ'@L�nR����Z6&bo�m ��wt��+�F�Pf�A�ڴ��ְ��3����{	 d�`�]Q��l
&KEUuc�m���1I��������"_9+i
��RQ�+W�񴖄�A�`���֤���=N�B�!�HfX;�	'A��$^��#u�XV�;�d�I�@s�_�~��S �~9*�0 @P7�c@ s~S�Eq!h�ں��V��ƆO�5E���YE2B���O�������Yt�D����{�U@T��O�Q������D�5f���	$PRd��#�f�R
vvփ`���vЌ��s�O/��������D�PY"
6��|S��犓4���n��M��לq��+��s�+{��ޛ죠�Zk��6<��`���|�	l-��~��b�N.T+��p�2���G�ѐ�������)B����z�Ƽ���{��==���9���o��xdh(�h-���z���)�x�0��5�@��Gi����ě��ճ��R	�v>��`�5���U�q��Z�L��㲳�452�У���7�W���l���1�)1K�t�p����г�v�#_b{�K��8`�/q�(����V��&*�������B��B@���������N1�z��gh.w��f�T��Ŷi�Q�k�7�����h�(��Y�`����s<����J���d���|@��43�����X��=����L��|�6=��N�����)�k��t��ژ�/�j��釷���=���+��v�593��c�V�gc�?�\�Z�E<7͝uY���9m�פ��w3?q�D�]6���Q�dL����Ȳ ����Vp,��i*�|�����\g�GB��>��#$�|W9��p|��ajfQ���˦6>�r{�L�ګ����:m�fM�*G)�<�,��/\��K!7zaT�V�m��?�����Ϗ~�{�n4�-��|��e����Y?]�I��k�~���ڢ��� ۙ�؂ ~��x�%� �󜂂���aє_0.JHD���,W�ZuRz]����R�z����1安�d?c���R�$�X3�ڇ��Q_j����)��a�iY���^��2�9�ll���M�~2ІbQݼ�pq�a�G�}g������Y�?����)�ܤ>�7h�ѾR�`|����?�	���g��SSs�l��ő����� G�ST��p��c~�!��}ח��>�Kc\==�%6b�:
	
����	8���A��de��+��������E��w�s��/xz_j;�`��k�G�����5{�Ah�m��FSC�e{{{�l0���dnXsx����� �G��;���}�z�����X�L�_s�$T �g:�xҪ�(e�$q�ݻ;F��e]hY������Y�O��w��41��~��
�h2����o�=��)�-�<���օ�*�u1:�5���'^{�U���q��?���ڕFM���:h"�����H��Ub�	��4v�}����xs���{�&&&f�xl.�j�	��j�gX�����I��V_ �<�<c�T~�D�؛��*���\�(zf�[��kjL��6s�����K��'~��JV�7�XTT���|SfVձǍb�O[ͫ�s��Nw�}M������Y�F��v2���R Է�A�)�I��}W�*'�[4!�w����kr�B�ٽ��?'�j��s�C��fע�d"CisZ���έQC�A�APC@�Tt�E�P�s�-�e��E�Pd���i�^��D�6�ne�����2)�Y���+3i�i���^�Y� Z'I<^=�ĕ����{�� �,]���ɑ�y����m���ҊQ��Q�	��;�?�m�xJk������A�p'������B����
���C"W;������vhf+��.:���<�GXO�>�P�,Cb3����[̖�:42����|�z�l��F��v�"g1����Soϝ ��㪚mw�\�-H��>��"�P�*�@D�d7�Lˢ�)U���`���&Aa��	�(9*`4��I2��\w񞊩-�t��SS�]8� �M`�˭}��u�E������\������P�L�H�,XZ�dR�)π;jh���s |)��`1祢���q�U�O�Pd�����Fv������� P��q�_�)�>?�S��w���]����uQ�Cd��@�|&ֽ��ւ�>A���D[��t���h�C���;� ��(Mc�f���9���s�v�0C�i($��"���Z���Bx7��LM[g��'�?z�8�Ď'ԑj�WvI��A��ѹ��vh�CI82�m�����sxO�t���;�űWe��S��=�ed��o���
�BS>YK�8���I y9���F# d�����EׄՕ�uu�~��^Ke4ǲ�T�V�	b�e!��cq�?'Ɏ��Lݨ8���k]{��u'�W���۴i��ֈ��0\&�����!�P�����W߱���H��ZA���`�kΪoY�7�W�����K%DbY�sX,��<mD_^(��]"���V���KB�m����)Et�ώq��t��Zw ��L7T���6ګL$��kLG�1�D�E
<�M�sF����8�a���l��$�v���e�����٧c�Opd2��.|^��S4��ݖ�*K!V��9�O����L�90��I�@��a��OU�Z��Ԍ�[6���@���[�"A����;��'Ꭳ�(���k/@����_�b�M)$BjW�9f��P�-戆��X����U�5:)�����q��}S1�z��A ��܂]�'����1ǃ �}E�\�y�d��\t�؉K�\��vu&���w_�<�h��9�WFZ�K0e%�C/(H�Нh�v�Ic��i��90�wј[�V,i�g��`��8	g$�z#p
�P�����Gw.����01�>�������df	�eފ�D/�������!pZ	�ES���lٲ�q?Nw����Y���	:Iw2l�'#C"�l�Hk5�Vs�
v>wdN��|�ޭ�#/���iѨh�0�ѬsR-S�¼�뇄mq��`r�#pO㱍ؾs�b%��3���9n2���a�?-AY�p�E���E����(ā���#���t"���ʕ�U�E���?u	�=���3�..��eD�"�*�m��������7΍<[*L� v  A�s|�;0�����A��]��<�v��>�?�u���B���_���AA~��i�,*�k��n���
�j;c�B��2~N�Q�����[9�B�m�߾y��A
{�3NW�8���<�@�{ٲeh�WoM<Yzc��oٺՂ���.�����:\ ��M��ُ|���"�? �ݿm]����F�֒��Ì85mm^��&�t��ǔY
.�YtH��XJL�����6�ؾ�<�<��=8��+R�T��E�٢g3���
'a?x�τ�����p����r�(*�?{�E��������cEJ^�?���p<~okh���b>Jz�TyKt�������������t%7�'�2b�*�ԃ9�Y�H�*��tFL�7�+̧�'t76
��c�i����o�D��b#�Q2�Aq#PƄ���?�����9���t��rX�_2��!��VA 3�f6��)LiQ�06X1�*�&U��0�ع��r=v�{Rg�E��_F�!ި���llx�`�0ќe��������B�[mwR2����%�Aɡ�3�]���ș���s#�%��'w����{���4kD��E�:��W�^5��[�bj��L���"/�7B���0ú��{���#;���~5��:��85�k'���M�Y���	9���kdD����c��+	���`���>������G,��Pߞ���j%�|p{�118���e_��b�t����;�e��sHjR�NGl ��F�:0�U�H/�e���]<�g]���c��E	Rė@e`�Z�g����}�7�\����zL0)�c��a�SIP�3V/�v�E0���IX�K�ڳ��8��}	9��ib��յ��X����Ìn�'����~~�e)��_>]���W�:���d�jhh�3�N�˽�2~ݰ�YӇ��U�L�ӎG��%�J&�t�}�ɼ3T�h��űXm�������Poو�M-k|�s()�'&�Jj������L�Z�
��n'S�g��T��GxC�FQ6i��ڰ��OI4D�L�L��;�h$����\�>S�um�=����98�/ҖBi��+�"���l�|�T�]�0��&�@�^A����C`I��G��&Ms�KRH�>>>�����6�L��FQ��G�v���
?/Y�m���|�-�� ���<Xz��g����]��������\���X"{JK8w�i�{b�lR���ӻs=�x\(�FwN(���>�G����������+��v8�� �̽�	j�\\m}Na�Z���@f�<�ߝ[<�C�x�ٵv���㕈�VM�'a��[�Js
��1�yE�r[ٵG �7�}�F@<�;���wW�Ԫ^?�����h��оEkn�������\-��=Fr7jbj������i�
���޽y���"�]5MC���!!�9z��x�i\��Z8,�(�v�V#/a�Ht�"�!|��&���kD>T��D���n5�;����������__����ib�����f��7�hF��y��:g��9����;�?^f�R�1�28S�o��[#}|r3k=�Fv��,T#����)�����D�k��\oܝ�y���ML���z0�zS9� �����.��sr��M�|��`$aT��j�(�%��U�WY�a@�P.f���iiiIȣ�zQ1��Z��\5	L�<j�TǬ %�����N��А����	Τ�`,!]���(� ?�iww�m��Ӂ��z�:9:{>�R)�G�n���S�0�m+V|v�ͥ� �l8{RmZ��� %�Ï~Y}��vvv�i�(s��lgk��Ï��zRw�$(��zy-Ȩ<ֻk߯R��t�ɧ��*oDoE���D��Ň2��.9��p��R���3�
-�& +Gɂ�8q���o���+�iZR���؊���Hf�n�~�Gj��O`������[�v��{i8r�\�=7�Ih�������`�>2�Zݼ���������������ݫo��a�z.l�OA�F5��p�4e\!�;����n�Ta�M��[����`eG6�e�x�.�e�5g��C�+E�GCJ�$f[1��������/���9�Z�Cw�Qa�=0�s��-�Ϲ�Z�$��̓_w��Y�=X���O�%@��Ȱ��U��^䠶�=�m��?%���7�%�+�u�u�Q�[�#e�����M���r����xl%k��[B|�Pzwz,������)h؜�j5�t�_�ez��,[�d�Ґ��sB�.Cw�l��<Z��A�x����j��l���V�'�H�'tS����J߰&F���>����j��Ǒ A!!>C�WA�#	+(��PH)u��Zs%�=oz][H��,K�շ:�DC��j���+�����P�]>�NTt��1���f���L�I���:�!�q���c�߻����ݏ���ǌ-�{dg�)7_a����[>���c]��~G��~V7����i�땛����ݮ�~1V��������8���>/�;���Pr��x���?�����Q6�ᛔEP��,6���ʕ+�"� ��+W�Jfs�\�S�ޏ��J{��TE�ф���^n�U�F��Up+���1�@��A���W�V*��Uz��H66{J��l�S����P�X�
�j�U�u���W]��͂�ܡ�c?�!��D�����``&��ZS=JyF�?���u{Dg9R,*첑��G�\-\�cy�P��ӥ���k�p��W�豕*C�\"����_�����4�H�92k�J%|<_����Y����̏@�;;9-�!-��8���H�p�n��s� �h��"x��b��)�����R��]��/���^E~ӽ�-^*_��ո M�;�����k_y��_x)�� Ӱ�)驆���R`Șęd��7L��FF^��B����n���\��>ۤ]_/s�.���`�/u����`�6���T)F6]hGNί�A�Dw�4�\�amn=�X��?T�P*�=��xR?,~
�[����1^�~M���A���ee=
		��|(��-J�<�M$[�{�m��(S�P�*B���x��*7HD
�"2�֭�
Ua3CB�ܔ�|}�zW\�;�+b�5p�h�C���?F�6 s��F�DYZ`�)���J�Q[@|��G���ć�@<P�qf񌅚���5���y��N;=�S?�Y�w�X�����F0�OS9S����z80����ߺ��䊉{O�v&�9�6�����l/��{��Fd��W�k� T"��|��j��Qg��Q����BE/��U���z��75�%���hJÏ��G�s��|���B1a+������&�~!�\;ea�]�@cz�/oՈ������,L���Y`[�.Z'�:aVatB=�� 5gL�Ő���3{����|��i�Klh�<8��<��i	�G���v�B입q1���Gl�4��
�uO���r��U>O;��M�8� n�rф@x%\vPұ����~��9%h�.��;)�����(Wg���5�e[}]e���@>�_	>tʭ��bdY�W�3+�U��<ָ����Q�׍�VU��Z˿΅#+ۄ:k�F���!��
������<L2�ǧP�^Rd�	� �D}��	Y�,s?��b"k�A/��jr�;)!�+;�WFF��5]]&=�t�Ǹ��L	�FY�L�F��3q��Η *l
��A}�?6u�^a��%n�H ̔�m�d�<���đ��/��i���-j`����o�#���Al�=F�qd�]*���L���yF�T44�޿��(!�����X�1ec�qj�bA���|6%��T�>�W�;�=���5�只�=+��.�V_"kH�*B�����榊�Ј�//��X,8^�������>�*V�Єc����\faii,�����ՋxuW��ps4NW�:�ޓ'7�[46
9��� k�\(k[T�Rٿ�H<�o�a0�	�Ugl��ܙ3�N�8��<����"�5r�¶� ��/6�};B��=��+x-^qcP����ң�B�#�?<kkn�������?
�G*w"2�t�X��ˠ��>���������C���)Zg疭[�><�
�+)i'��FG��)���a^�n��=�T3�3�)�`�8��ӱn��`9	�|\CU�nmd����?A��̗d�~צ��#Ќ��es����,s]4;^�W�nw��"�\�|���0��}��'��@oO(�*GW�C���N��1�����u��3	���Nz���Ɠ��[6����q��ǟ�v{���5�~����,��4X��W��z�O�y
��������aG�x|�FP?q���߉�ؘ7J12�7�86G=3��U��v\�r��d`����o�'	�"A!���5h�W>��[�kD���i�_B�B7՟O��5岹��I��K@^���OL&���;z��8H��C��#�<�63a�=�ן�)y�X�FDTDd$OL�T��iZ�)c 7r�q�vu���n�C��nU*�a��T��	�a!1�R{SK����z�;���i�� 	\�7�<�+�6\�@P� �,Q]���}rٲeZ=�DZ:� �X�\���T�y�0J@��ykW4�\U�Z K�<sP""�)��S���8�V��hS��|{h:�Dς���"=�=Ou�� ���oyto G�\��҃kK�^qA��~���Ր�o�<,LIY9E8Y����F4��@iiiF��'�b�U&��у��S61b��WܴiJC?2|�׾6��Z~�0Ӵ��!t�}*�v��a�m�㑂 ���ua ]ET����.�0�0����_؊xVC{��p��d�k�=`���gE��sF�ج	���3�ŋǆ�?��?J�zZF!����9M�L��k?0u��`��vz,yu��@"��o�v�P2fcK�>�c��+���?�tt!S,n&H������q�q>�*��8�S�-��~4�hm�Q�-ׄp�j"��c�f�K���R��h99𙦦��H@����Yr5�65��(��?T�G���H�F.�oס2�iZþ�j� (����a)nD�#F'7r$(iw�,��63��Ԧ�t��~5��W�Ǿ�%Տ56�y����Ct���v�<2'�oe��PQ�m<�`3|��Y��P@f9�	cڝ�����p�ʦz��^�.]������������� ��i@�L(� �4Ѐ�]��c�(��v�A���;Je���p���7�f!R��x���ߧ�V*�Q}�nK�יW�N��m�Ꙉ�x7\��v�:�F[��E���΄�<�-�?fW�ôF��Oi�
�O"ӂQ����g b��<2��H�Y�rYF�<��%St���[����~�5ˣjo�qg��u	bj����:�Y�,'3P�~���⍥3'Z����Rg��}W ���U����3|RQ��cO� �������kaM,�ڬw�ܷ�nh�E����\S���R2�:�ڲ`A�Xm1s�\]S#9�/l�A��w�--�as���xۉ�s�g�̔c0�l���2֛�s�.
�{��7cT+}���4��#�Ϭ��@2rr ���^^����GN���"W���>��ބφo��/y�-H��Xw��k�{zf&��ݵ��ɀ$3h"iMM��'��(���	����iIXOYo�.�VC�X�ӂWALneae�#l�3�
��Z������+}��>n�>�*ǟTг���yP=�zU��	 {�����ۡ�^N&��4D$�l����ۛ��{֛H�|�K�Qb]���=�NBW��d��#�7V���֬`$�y6������	b5o��	�{$cdd�6�u1�:����g����r~�[��5������C��ZX��BW_�.����O�uQ�A@<'�E�l�"��#�Q�MM�Z�{�"��
�X.���8�"Ps�Ǣ�����>/05!�=���xw����K4�y�Y��|wWvGQ�6�8�*q����*�AN���>����[���+o�~&<%=�>�� H/���ax��wϠ��c!�z��8/e�_<w�[����Xw�0n�<���P$z�@�~hQ�iݠ,��������C)����a"����Ph�m{'���u�>�+5��N�Я���k���`HXi�_|)㦮\A5�p�)�dQ��`{���ul&氖�(�I��ԋ��wD�*�څ�\C	N����(e���F#c7�0�a}@$���\����չ��5��#ӊZXFd-j���*��׬��� �!0i��:kk�{9g3���3�3�/�
<�R�Kn�ttw~I���k+�7O�wRB���t�u�b���7�˓��O�=�y�֧QQk@ZgX�K��2>�a�,�Yx�v���rFj���{�,�!���L�	��dȻ�4�-7JΠ���+���gPϼT����jm�񎁖l�V&3[�P������$G��᫬I�H�z�s���t3���ܠhR��ЧvJ������������1��c��b.k^oQ�/�eHW�-�����p7��ş��Vr�l�ap�ΰ��R"K�a >���}NT�2Z#e6#�[�ʍ�
\����·�)�0�H�}��=�|����uu�Äc�������߮�M�!x�1��I��St�m^���^c����Hw��=�|�$&�gcd�}]�b�R0F���P�&V�^.�oi�l�xOϙ��[H�ڈ$� c��p6��"�����[�,��3��wt2���s	K�rr��ֶ��*�q^�g�D����X�������h����n��:͙�UA�F�vك���g1����)�����#���1|���7._T���� m�ɺ��%[Q�f8.`��X�"Z��Wy�&d`��(y,A��RXf�ۻGBY�<��I���*�e_�n����Z	Ԋ������N����ц����I�km�q\Hc�k�Ng�L��ק�nǠ��!����D��(iv�4��9��p��+RS����Z7Ř�b9�1c��3/%��Ha�_3��TW�qvq`/�ş�(�X+D��(F��g&�WI;��K��їU�E�T780c�ɀ������c(�c�w�ޛ��1�?5u�H�1�e��!6Z�J����\L�5����3�+n���4�ĝ����a��j0X�x%�^��d�@l��-~B?*e�,��*�U��~&�m@�) �`�	|!.$��y/n!�?{^yWm׬D���G��!)?K�@�H�l��Y,��o����2�!�=\*a�o��K�m����
��80(��)3d�E2|�<�v��R4�4�E$nIe7��ԪE���aap�R��'�2��7CWQ́���H�rR���Z�}�r:�2�UWY��:���9)ݳ�x��z�8rv�OO�'�eǕ�� ��o��F�O�X��P���eS�ebcų�ḅ0&�O���D*�/��,�e:)�*c�b�_�?c8�����很�0�c6·��}Z����6T|4G��'���'�[t3w���t���nb�e��(T@����ĺ���&� �k'>��q�-�{�~����JKC223wĞV�:�f�����YW��*' P>cf82�/wH��}��:��.{7_%�98���}���F`b##�C?D��%%�jV[[�TX+��m{���罌묽�2�岹��x�օ��������'{�nYq(��x2�0�������~���1�fpS���S1�ģb�1��u�6� ��5�O���Z�Ldo�&{��3e�s�L^���t��4[�Xo/*�sS	�b`\���=HYʹp��[��0�����=��I�Ѹ����Ս=�����h���R��̩9�q��MZA"t��xTE��N�.�^�dL����_TTܼ�;(��� �|q� r,a�����J�@'�����G�4D�vFj��w���װ���<�4�Ϣ���(ʬ�<��X=�"Z�Vn�,��Iw�Ce��k¹�=8|��K]�qͣ{�%�_�Nʉ�>W���`sK&��:Tcw�� ��)8�q�v[|S.�m���%�R}u>�k�<�1��~] w�u��l}��?�W�8����4���N�؍Ub��K�g���L����Q�a]e?��T�ѻicy���ޘ�'�����"� rÂb4��7�����6����32.nr�d�$p���ܦ,u��-�U�3�+�6�H+� ��m0�жg9`�$?� ��lt�c��A�[z���yѣ�5�g��O�~�%�-<��oz��m2�����|t|��X�
�!��]qc8i�0P����ɼ��ST�\54��,|�$�ӄ==��O�f5ٟ,أ���ד��a�;Z��Ic��n��.l�e3��	)p�բ�W���eOk'�F#��,���������>w�p0�D\�ڮ�FKsʲ�3%(���շ��m�R"D�e�6LC����V��JUB�d=�bG�������rj�حC~�p��	�+4I��VٶƉu��^�����4�oa��`�~7##vg+���~8����jQ���3'��z�E�-���tS�+D�4�hF�N�J
j�WG�{�2��@B�����K�֊*�N.T5"�&3�P��ֹ���º�^r���Q_�����^���p�F`�Q��h#o�l�c�����F'�J�գ�����`���I�*�[yG���C&��
�ި�f��/����E,�"]qk$����G��'��_�>���c�	v����J�j|Mv���K���gN���u��^?��:����Ù�/��;gb��eʄn�Y�x��)�Sxō{�σ�7Z���a٪1���j{!N�̨ؗ��,�2% �״�<�v�`@d���%�z��d�\��...9C��V��q`��劆���A|��Ηv�u�����Ov]iq�+ݹ��a��_�o��>��XS�_����^��۠v�m!%9j� _;NT��ܬ]��������X��QuQQ��_,��QO��	����<G+�8a���C�|f���#�Hr'��q6���4�yy{'�e�v�?4A��s-�G%!g��і�t��Q�`d�
����[E���	)�^U��<��|��,��n8 �c����Q����Saa�E�!���.ySc۱J��O���ٔn�S��0��z�7�
Ƨ&�X.-گ4qP�ǫou�X��r���\3A��x}���X�c1>�EF�R�g_������O��<3j�FR���� _�{��q�dQ�O�?�8�Q�o
�������>��}k�\!0��h!!Lv��Կ���K���>|���k�����i'y�9Kc���Rc�l�%�f]��*�U�J&�iɐ��3�2�L��b嗇��d!g������o+�]���q�H��ӕ\q�u����eGjzO�����u�6C�z_��Lu�ڎ�h���E���{��P��������� b`��T��#l�|\�o7�܎��M�4'��� #���,��f$}C�,m��u}�f�1^��_�L��d�����B{��b���A���u��x65��k��Lf�@p/��0��N�1�|�z�����e��|�T4��%"����B�5��1������7���>�?�+��)K9~K��\�{�BO�Æ�zSO��b3'Ҍ���*��h`���{qfM������ƌE]����W��d�=X�cX�2��]�{�B�%��%7�j�>��-��G���Ӄgm�4�"��S*4V�7�}���j@"��R�cI�ѯN?|�&��
���%#ֶ9K��/�y�I�e�R�0		v�:XC(6圜5gk%���[��%�f����Vw�	������i ֖P�Y<�,�muR��]9x(\�gp=d����@��}�iZ�t	��3`��J�Ȍ`J����;�LE�?����ys1�Q���>V��8��|wG5>xB+�?���Io�T>�ZV:�Y
xLW����w�:�O�wyiX4_��vC"T�Tۻ쪌���.q�ҳ'S��|��JWVc!�Q�5�H�tq�w����s���5����~Ee�Y��[]��ǉ+d��Ev"�'G�g��	�;5aY�߅���dt�F$�r:4�/���;���ݢ;;�(�,F��"�!����7]��9�(������_NS~���},y�T������ǃ����yMX`�_�0S�L�U�����(Pa�����c��,�ة!^9��&�`�1�����/��'�g���e��?|8|�����b��	3���in��H�	���S��~�|�e�o�-��Fm�ʓŹ�9�Ҋq���{���$�}*�\��^<X��<�R���Mg]�}�7$(���"��<P�mg���4@e�O���q�'�xlNၐ�b4
�
P�,�KA(�
xD�3 d��n$ͣ��f��^O��x	�n�D��Rv�� !���>�nz���T�����/��࿶��P�A��æ�a������[�n#{��N�~h/���R�c�蛶~�D�h�X�'���Ѿ(¬��=��]�1G����f�Ƕ�fX�g���6����R��BR�lӹ���I#�Aesj�P��w���ſ���{�t'4����Ji�\B���A�S����_�	&丣�#s����`�0���3ݕ�B�5����s���/��
��"��S�]5��1�ff�SG��Wڟcö/m�'���5��PKk��$V'd�� .v���gf���j�pǻ��ؾ���t��yp5�����$tR	���wcc0�ߡ�������~rq���)jq�m��.`	[���=�?�Ú�.�Qm�zp�&��E>ǯ��K�XYjE�a���2���90����a�t�*����\�B��t����>)?����# ��a��DA��T��H���~���X�wg��wϯ�S��
H7����b�w.ޚk��t�E"���!D�����iB�ߝckc��8��֔`=MyPz�4��P�%�Q��hk[�gt��F�0��2�/j�޸�6x��K��a�9I�mF��a���L��3�r�n6�%ޱو�M�G�8�Rf�HLK����#�\4ٳi{-��'^5�Ò�8%D7 ˁ�����=@����9�b(���I�{S0Ճ���.�
�ѹ9��Zj���
t��fj0�V���nc  h��u�Z��
2�B����<>��᠀�jk���5]�R���� ���	G��Z,��+m�4[��n���6��3dHU�F%"��Y?{~���}��u���%t\�����R?��- ز\��� ��z���7~�q��i�6�w#��Nf��I>k�B�����{8$�%�1�����Y�����\��^�Fb0����䊤��q~=�s���篴�a���8_q�#�x�.v�(kW�M%b�pv!z��� �6�/J��R�H�i1�����:����F�r)D�&����Q:�F$�7��i��ʁiժ�Y|j~��Φ"���Y�L�������W^=�1��F-p߇����)�2M������!���T�o����Q�89�p@�8hxٹ�3��A�8�*R���F���ǁ�	�)������<Bf-�g���us�y�YO8O.�o�o�'���i��1��.>e���Lc�{f觚����ޱ�l$�����F�P��	|���#cS׎�F @@Ė��Ra�b$��֡�b)#JD���1\-�M_=��(�j�Ţ^𣡫���T�F{"Z+�~[�Q�Y[n=�wVHf�J7Ex�P��O �<6�~�$;������� O�����m������|0��ݽz��7��<�,�Ctől�:+m��#�9���Hd'�� �D+���� ̃���+֞(d�2��*�#�R��^�V��8B>���6����l����bΖn��N�%�M��|����49�m��r�ht�/�6�]�?�r���t�D���7}h�=\*e'[~�G���3JEYN�]�iq�0������ke��L��wI�?rr-k�]2ٷX~*�tKK�����x�H�v���<������{���mm�}-i�&���P���JcX}iQ�������ّ�����"G-dc�(�avS�bsT� ���yLT��dH	+�H��?־���:�I�([��Be�V�M1R��%d�F�PI8�%Ĥ���!�Thlcd��L�1����9:�sN}����^����>����g���}Gl�o#�kG��!�,+r�*[	|�q��l����}��[��B��[\i������L���>�7W��tGFs'4֊�P���w���H��j1s���5 @�ïJ�ύk�e�[����%�rO���	�?"�� ��)o����@��!?�[�(1���AK]�G³���/�aڃk]��hF>XL%Wj�}��߈��@ �-�t�@������q	�L��}���hpD��=h���GOkW{�3���b�|��E8�-GC�܏z�Lbx�i�6�����?�ʜgo��9v���n�\��/qR��&8��J�Q��Ŏ��'F;��!�x2.�X����p�U�s���L3�:�~��T�r`�<3�G;�H�{�W�Q*��y Y3g�@�AOˉ:����.~g��Z���+��{�5NG�F6��]�}��p�aΖfgF��=o(r��ڷ�T �����
b>�8"�~��2�/u��(>v�W �W==zT�!z�|���q\�W�����1�H4���g��5��ʻ�H��w�K��Ɉ 3y���'�G��������FB&�j�a��M�v��o������,n���E�U]C�`�+{��@s�U����{��;=1�Ӣ�筇��r��6VAA]WWRff�9_ߌ���d??*�qЁ�į�貚O��.�jc�6k���e���W��&��B�)�?M������9�����E�'���R�b2l�����{Dt9��7R���H�1��Wٛ�ȆZ�C�ej�}2d:`��C��&Vۘ�8�f�	�4�2���H���Үz��e��Q�C��퓟)T�ȦP�� m�D(I8jOk�����X�4���-HlA��"M��o��z�������W��{2u@
j��_�M�H���;�MS��WЍ��(E�^�F��MȦ��k8�d�����N������E�B�j �U��E��8��������EG3��7���I~{
�|��ߟ�ݑPĐ����2R1��p_Q�g�������������W�v�LI�{���d��Ŵ�Ȍ�/?$��OR7K�m�����|�H��L�lk�D�M#���Qdp1{�];r�����-��+���t��K��)�wz�XO�tTa�*6h���+C�-_y��W�=�^�U����~kJs�D��5:r$P���9%��1�?N��a�]�BDu�
E���Ƥl������V��Y�)r��E�Q�j4�""R��Қ�:�����BM�I1�pJ��_����O�hf?��j�(QzN]bRc���cy���"
<@�Ow$D�j�`)� ���C��	ȿ&n�-�$��Z$1�y:�P�ߒ���?HE|�DEY�k"[{�	eK[����~�G�L4���pcݜ	���º��G}�� �@��e=��O����s������|i���t64���p�G3"@_��<���CE���k�\��Nd�^����1��v����	nu��b�c;J�93��;��;�_�I��c�}���f`A;��k��0��{�r���^��.1V��e3,%�Q��m�5[Bv6J(� �nnh��64�Pzgk�����qVd���Bi��z�m�w&[<U�NCkv���^{|4#]9��x��kq��6d�����t������� �~������ާH�+�BF�3����9r"��9�ܑ���$3�\3��-!���+�)-7�ܔ���,�bE*K�ر��zL��w�����O������P��<��k=��<���ϵ���ч�S[
���a��?m�Q���[Ae��">��u����'Ldә�7�Z�_%~bf=��C��x����.l*y�%t)���K���g���vH�~;��"	ܦ�TB3�����9`����2�a�PG3]5���e��x�6v)
�W!'Tg5د5T��	XBt����13|�uc�i�p!����g�	�E�Ϙ���o�3�Y4&�Hk_�h����NY���+�d��E�F�tRʜV��Yd���p��n�	=[���h��i��w'��� 
	�c��n��0�;u��n�˽��{�E���1pIQ���Ǽ�z�Zr��!2ǯ�/�~7�h>�C+9a9�l��m�Xow{�3�Rl�Wa쬋�y�q�)�ܬ���@��*����ޓ���}I�ZdH�"xz�O�<���̜�� �O��H.E�c���Ce�Y�c��h?�vp;Oǆ3�C���Y�΀��r_F����Z�_�%5��Un5��Y2����8�l�',qy�����Bm������AO��n�l�~�K���:����Q������Ȣ�_w���ņ�|=����5���=\h�[�ѵA�0�ޝ���ET��Ӈ��(#�Mx H�"ƙܣ��c���LP�_�i�t���n�=�5�4K:;����D
����_q;��J�s؎֝�!CC�@�^�A�3@=�u5?
aLU|�f�A�^���:>��hs{�;	Th�p������}������B��-B{E X�y�N��5-��ݍ
�S,��r���"�~J���F��c��m`A�
k�c�������k��ұ��O�q��F��B����pq�=�C�m�.��>�@ΜƖsQ�q�����oL��.c�p��J�HM�u���f����t�?��<q��mT~��+��������%n�sr��c��qں��I�C3��	r�Tt� �#�_�%����IqT�#z�ڞS8�7������0gp�I�aeX�O|c�nI
ucи����#�W0p���۾s��)v�G@��>r�[����B� �&:���F����?W��x/?�s���I]M迕�Î~�j��i�����ަ4���V��N�t^R����UJh��6��%r:���kr4�<� ���l�C=�p�o񴁦v՗M'����w��c��T��^��]D�����}�]X�\�����me��Q�x��|��ٍ�a��?�)�NOY�
1���ſ���lÐE��5�A��x�6��མRk�#��$���A��k�!5�-5|w�]��y��[(�Y٠��X�-��s.�h0:R�f���@�~$eZ�/�$��1 ��*�P�[B�5�iʃ�Z^��>�2�XۡS����H���[@��dx���KS͋��LS��Jz��r�4l�O�.����
i�K��y;�v~c�R���{���ކ84��rh� �#������b�`ъ��u����K��/4S������L<z�-:ߣ�"��h�l�őHݞ'�a5 ���"+7�@+������-���l1[���:�Pz}xq����^�Ø[�
�e�yS�u����K��'	!ٝf�-n.���]��/����?��:&�a�H��WY�Л_Z3��m`�Ur��8���S�T�֐��LV�0����.��Ŧ��yI��GJ�.�kGS]��L�%���]bA�z�����[�q\j�_�A��s����*MW��w������.S;��''SД�|�\�yϘ�s0���߳�r�=�y@�N6ɍ�-��b��çݟ4;�6�R	{qć����Т��&~f���⣺��C���{���@�ǻ��#ã&��b*mp��8�;I\���Uר*g�"�W��xˤ�>4ٰ�9�x�	o�+Cb>K�	��o��u���S��ȶ	{����7qLm���z=����A�bB���,6���
�w$쭰�fZZ�����h��(�E�^�g���'����@v���FؾCiʴ��L�N/�ej�*��r~8{�7��J)���`�8���'A���,N�e�M~0ew#x������\�e�+̡>�����]�i�=���B���fm��U6��Z�r"�F� �}��h���ʵk=P��G���{��Z �S��1=�X��c��L�u�k�Z�d�ISEt~]���I��Ǖ�PD�e�M�r�,�o���uq���ʒAST^��kRn����u�����ǐNB��t��ǂ�շM��㹃��@ ���t �Z�����S����E>������#�QB%Zh�ɭ!�ԧ������n�\q���Y�JS�Ԟ�VjOx�<3{PӁߛ�~n�^�'��		T�D�JG���?ݔ��r��Y���y�1����"���3KZ(��2y��c^�8��B����&:��Z�U˃�i#�`��3�cj��B絸A���ʶ�[8���<͝)�F)�[�z�4�^x�]
�O����%��n[ҁH'�#X��EtlUk[L�r]�1�L�R�]ヽi�a����|�����^�Ǉ=�����f���;ǆE���"/������O��"w�*�}�@�� i����8B����,NDsg��ʹ&b��2�e}Tơ�0��y�V'�0�$S��Fx9{���z脘O�;�u�Bd��k�{�s�Hő�a�\���lߙ۟1x�W���X���p��,��e�Y���-�6t7}~��?'d�1Hȱ��%��4�0��Se���3��cb	��CV�QѬA�W�詞Iq�<!1�w�:.��N��r�b�c����ǘ,�?��A��$P�x��iY�L�ܣ<cS@�����FɃ�}t,����߲y4fxt+�v� r"��I�f˙�K�3Ԥ�����#埒s�xg*V�n���o�J��Ux��pm���x��[��2���\�ݡ�nx�ṉY�yx��!�,^v��Y�G�l�RZ���]��� ��t�U���2����Vsd����Ҩs$��e�+�~�%�W��gf/r �fM+@�DA��uE�_Y�!�85A��ٿ�"2�cH���$(šw��XX�Q�̼��O�d������n�~�Fz��NSe�
�������Q�W3[J<>�p\��EY0SBs���Q6x��f:���t�_�M��U|�P�Q��s,�8G�kM�:���2P�e��pU�O3^�@8�_@D
�����F5��J�3�x�1��N���߸�������K�l<���^E2t�dh��jxt���C3��jRl��>�p������0M�`:-��5�����$#�X��C��:�*a�At�B�В��,�R�Y��n� o@��0��: 	���r������2�-�;��k��
�U��o����}\?�S��dW�Qe9����F��byӳ��kyn~������=#�y�N�66������[�!ҧ�����Igyw�>�@Ǧ7�'7�G���8VZ�x*��J3Q�_s�z�?L��h�1�������ݯg��	Ü|�.E�n?�|^{"/0�u`��B�����a���f��bb��&ܻ>d�8���5H�?}�j��t�Ķ��O)�]�����'������n��l��%-��w��D�����&O^}�e�uw��N1y��=*倯��� MR8��Z�o���,�%��"A��5���m�(������(3ձE����"/�sWG�l���wOҚi�P]^GNőh����"EЄ�R�ޔ 	~窈������Q����o7�aD�{�5o�(0�RnN�+S,u��p��_[�n���H�::��=qf�3����x�X>hMxo���^���@��(��y��tl�I��|��3�����uY_>)�F�f}�I����z�Hcb^p���߉r�&IX�6��ߨDW#�d���i���{�~,�޷���!�kX]U��߇%v/qƂݮ�$��]z�}"�$�R�"3҄��A����z�����_�Jy���H!z ��Lċػ,�?7��s�ʽ����iԄA�(��Uq��r��o�C�7GW�9��b� �g�:.e`�=X�nySD7Ŧ{�()F��Z2t-g�t�м���ن�0&ख<^1��S0>:��kS^Z�����p�4
��䷹0��
�5~�#j7ڔL���ʾ��Y�K��F�����À��(�f������b���źa����>7�� ��;@���V�Y��b"}�6;�7��<��S)����$���,���P,�*��6�Ot@�Ć#��6�i�k��9�J �dm�����U�1Ƣ�¥��xn����)��O�$����#c��C���ͣ� �ߝ�o�*|"���vV���&�di
���-m���Ͳ�uM��(�V|(W�L3N�c�h��;�Xވ��Q޼<�Su��b�$)��o�k,s��1JT��$�r�$�^p����[ȯo�]8�֑�}n/,�"����F{�9���9擟�ڦ[�����?��^zGZ�G��Ŭ8<Ju3�i���	}�xS��~��z�`�=���G�$������儨�lK����{���}4��r�jyS��,� y�A�D8��R���C6=�_��?��y���2�o�j�[���okDW%פ� ]�~�OF����܋��ˍ���$��	���3V=&D�LNS��xY�y��i�
N.�3	������@�m?���#G���j
������+���>R�?���%��EDT?��0�Q�p2�b�4����6zQ"���{ă��:@��W�$@�N��=Z�D�� ����dO����Ȧ�+��7L~����=5�����z��������������S*a��|^�����J���2�W�ժO���,�	Z�@��@z&�� �/sjx�,v�!��dzF������7��k#�S��W�.h@~���!����ݻ�s.p���>�H%r�}��ľl�	r��9`Âᔜ�?�!�x���S�L�&�E��:�ҕ� �)��g�����j�vaѼ����~�#)aA^&;��� 7[O&�c� S��N��_:�F�H���1;[�U�haf�)OtR[����u��Z��KKk�?���ڍ��*H�qX�k[���P#$|�)�;ChF�lK�W�N���%Ta����;�F�x9	��G����f+*"��9�����D����q�'�:�ޱ4�}`wݩ��Gy����r�	�]��C@l�g�x��!$�N��}�ս�HQ?��|M�g�[�u0�;»����E���}����S���<��t=�4��w�b-*Z���S8�y�!�SV!_(p'8�˼U���N{U��e֟ �R��qj��2Op�|V���j��֪���@~+l���_��v���Q�[�����zg�����;^��_*B��!�(�Y����K;ț���0p]|���l,��v��=���Y�i�HhvУ�T6�<bGbs��tю�Aw�g���$8e�-�eAd5 w^I⚑}�ұ�@;Q+������6
pC������ _��Ci8xZjW��(��I���ԃvy"��'V��q_���"){ix��{v��(��9�5~4#���5��=qG�z,	�k�N]��h%R2�>,{ҜQ�t(����}s�T��6; =b��N������Q-T2�C�,�a�A�j���^yD���|D��xa+���SS�A�� ���C!őV���������Z|b�jtu���9�� ōb\3��E����� �
���2(H${��ܔ/cj�)RY�������t�{	�iy�n�O6�V\����$x�7=�?�4)rN�w�T-b����G�����M �U����+�Yt,��	��:!�RI��" c��^�V�Pҟhm��z�̎���#���@@�oa亵��K���˪���a��Y��3.%BPTT�;-��$�DU>%$�{�z�H�'�.��* Q=F�����[����U��|\ś�����c�vO"�������=@��%3.{�4|���D����I1�1��VE+|�Y�ty�
\����ݞP�����e���@���O�n������y�c�	�ҍf0�/����e�^���*���O噁|������}��צ7�a1��}��Em��Lϟ�)�
���o�Z@�ˈxy�xYc� ����(��a^���e���
��F Nʾ!f�r�1֐il�wz�1�tL�1u�K�:jEE GPQ�����M|3q��vb��F�2�o88ȏ�_״��/R���)U�f�V(�uh@ �4ʬ��ܲ<繫��+��b��l���\HV�n&&��y�j�*ͬ�z�\ߏ��X��\�,q��.7����;ʿ K�=�	��U�[��㦾�X��ѳXb�Z�s�;g�g��9m~�6(V������8�,�U�(�q�H��v"��n�>�,x1������Ȣ�ڴD�'����Q��I��F�ꜜF��f��4� ��a�!�_���>� ��������M��Z���"����
[ʾ��	>��6�y�Ǆ?������n��<���^*�U;)E���t0�������s�� .o���/�Y�0�I�gُ>�H�&�/@)}���~���ԃ�AjZ <�^I�m'�l�Wal>E!�a�Շ��i�����0���m4��_�8��Ҡ��-�coSS@;��X��TL�+��{tC��\�A�c������E ��]�hT�:D�>D��q]�����L�ŕ�2ԣ�i��#g�D�9�wۑB��LfN�����4��s��|n@��`�6��\�t�Z�o� r.�bV����ѿH��"bLR͋\e�V��<8��'�xs��	�i��Kvu��=*�ʮ�a�"�� ��Z-��嵉�[�Wt��R�5��V�.q�˵ݓ��4m|��͔I�1k�K7�H�� $���),	�Q�v����<#'8�~�8�ځ�{z�/땓ڝ�8�AqD��X�^!3e�|�88�r�2t��?N*�ƃ�θ۶W�N��er�T�����b�I�s"ʔV�I;b��s�7(F�n#ޣ�E:j��ѻ�6akʜ;=[�i�����a{#)���� P�^m���QU{��r@�����70����y�� ��`��S�
{�������{�3�r��z�ǿ=���ę�,��N�,���*�����
���}p�.�[��k��t���m~����'�2�_�]M�Ry#Q�#z��tY��m��D���r"4m�������H[K"i�F�����6���)�.sܿ�8��7����,�����GF3����c���J�բ�A���c��Z����)�w�e�Deg;�?sxV:������縃�[�L|���{b]���h��P����I�bq��B�H����(�+M��:�.U_�Q���\���+�70���L�r�@z� u�Ez}��B���P�~�a��kP�����6�8�ɏ�#�v�љ�=
1Y'3��;"���(<������������KzA{��V�g�䪪_�tw��#��b�;�����\��t���]�j�D}�啦�G�0�5v����$�j���F�ž��Y���,th���$��T����m���ԃ17w(.< �{�=���:�q�]M�D��ꨏ6ub�%�����"S
���j3!���~b?�5���v���jttK�I��e_[���#})ϔ���nw��Ȩ۪���d@��2ǵ�F�r���(fY@���P�_kbS��IJ���x祙��xN��%����{W��(��YY{s�޶��/��0��u�脙'���2^��d��i�cV�(m�#1Yk���=�/��+�����F��4���c�q��̢�}���h�h��iӲ�A9;6i��G�5�j�������_��F�7y`���#�|�_��j�`#��2��԰TNX��^���j�(UK_;.��չQw�,\t�\�X�E�r��v����o��	K�].s��-՟��e!��(��|;�Y���|�T�l\��xa{~o�ت��sr�,�Đ��ٕ���(D6+^���_�`��E��s�W�1�L ��Z�0+�FG�K	���f#�ղׂ�^m��eGܲ�W0�y��_m�my.�XV����899�S��r�����{29o����^�̙3tB�S.��ƫV�+��AR.�B���p�u��i����C��䌮�R�*�}�|��*��)�jīP!X��_�^R����\��4CW>V��ܜ�r��j�˝��j#�S弰�A�~~m)>A]y�Q�Il�#$�x+@�~��qn������{}����F=�6$��F	��ɽ{ ���ՂG3���w?j���ֲ@�n�c�+6���7��B���C�kciO7~TS�#�$X'A�{�7@8;['�L���V��˾ɯ��V>muu��~�ba��6��d�I����#�5�+;$��K�@�>����yR�Po��T͚iqv����#��}.�w'Z��Mlg�"�Y���I�O(uH3K�[qt ײ���ώ+5�z�Ev��RGM�Ϫj�8�O�����ά�]�]�?Z��AG�ֻ�&o�������[�֍9�AW�����ZX8�a�`|U�H��t"u��a=��]��0'GW&���G
�b?��Cph'V3��=��8�w�:�;=o���`\������
����Q�u��j���uv.�ek3G/�X�FJLl�)��^˞��=~����R����� �k���-��fYVW²��x�,,�؛o�q(�h���7ԻK^�J��zrZkoH���2������	R�fs?g0�3�T�/ů�~o�N��7z���q�I���}�k��]�[׉ޝm�"���Ym���b������.z�׾w�j�<�Z�!���X����3�
5��Վ���UoGoP*���m�9��Xk����h��d����k.�A%��=J��Պ+<<`�o��X8pU\P�S��v�E�����U��(���P�h��յIѶ�������ژ��DL֙��e��2�^�lng�"�ʑ	���<
�s�7�|'�b� ��b*[��-���  �n� 3F���ͅ������W���oںUn�"|t�s�ܣ]�4������dϻ�CË��)�3��2U-�!��w�4S>r$�ßg?JP2yi^�dX�8�2s�m
��R<���`_j����/2le쥑��U�M�����#rs�"I4k�Ҳ�ݝD�ݜ7�����$�9��jR���Ȉ#��V��"���Z8���B�
�:�H��)���Ü&��Wn�_Yn�&8�����f�n$�VVm��}dӐ>���,������T���M:���������
@�o ޸.U�VAcҏQ.��P��LVY.xZ5��O)�)lzw#���].�h̕�Pz/y=py�&J��R��5�'D�����(+EH�=tݑ������Ղ�<�P@{�"X����=
�(�mT|��(���Xa����9��iP�q���Rk~y�vHG�L?��lZuV�/�/4�!�����g"����Z��XuG~���^[)w�/6wCϰ;�u4��!yه|G�gE��$�N�z�?�
�3��" '�
e��O��^�)�.R�rW�[o��a}���s5B��*@��z|�Vz�͑���7ʭ8am�i��ژJ �#E���rʴ�3�1Ue9�#�
E?�X�������Ԛ����m�X�s��q߾eY�.F�I��l�Qά/L�F�\�Ƹ�0`3� �J��E�]"�c��/^dV�Kv��\�ማ���3�ގ��?�w"�Xơ��@�QA�Y�n7�0�ی��t���\Z��.zBu�m��^ǧ] Ӏ���s�(�XD���Œhj�&���Q����ON��1`-�KJ�'�;���k�H)�#�q�n�Oȓ����1��.�ۇ4I�m	�J��݃���=�v �t��w89����G���@lĂ��dY�?%�4���t�͡oF_B	7���v�z�l����4)R��u2�E����[���0h:�uߖ�2�:���.��;U��Olk�j��8T۸��d�K���.7�������V"e���W(�5�Z����H�u¥�앰�'��L���QZ�����c��jhh(�
�*�P��Sz�G_�����e�Mo��|�Q����z~%���H1��H���v#����U��G���?+T�G �� J��B��mK��IWU�d F
�RBj�p�W$<����׮�Q<0�t��߲�����&C}����=��˃�&b�T�D�We�}��-��ԋN2/��3<b	+���ZJ��_f�A�λ�K�䏆�`"��΢�C�Ƕx��(�^6=Q�2,#jB>Y*��b�կ	��e�H���Bl6�o���N ��:�mw��M!�{}�P�@�����U4C�G9�L�Z��������E�V�����>r�D�l����?Pԗ�򬁏���ړ�7RL_B#<g3By�E�-u���4r*�����hrbj�	����k!���(�X�fO6Q�����9j����2��:�nM�T��"eK����mՖ
���Q����^~�)��+�!�����>s�̋�)ߕ��w:�УuS�����x.O�G�m���Ej��Z�Q�=c�LhFV��=s�#Y`YH���8�����g�����@ho\�I��^w*�ȗیOPU�����}&�@G�0mQn:~��a����� p�j<���ٛ��������s�yf$)6e��0';�}���I�o�f.^v�D�ӕ6 ��H�Z?~��b��l�6_N*>�n}��`H����/��4s�xlC��5Umi���d.�s�
F��l����92' ��!�$��	5�����B�����iQ
�^�_�?�G1Έ����+���=�7 �.�qÏ�~�d����Y{ծS�i8]�z�Y�"�t���q:�{�bl������O�)܍���mmT��EO���k�MA�"R��,w�%,ُ������&���e��/�<c���	�y�ѸuO3�Uʸ��N|��ɉ���K�H�rYf����9���z>���>��u��ٹ�ྒٜ3��9|A���I���x¤.��/�t;��m��-!`UVCE�f㪨�J�kH��.3b}N^����+G�5��8�B��r*ɤ=��yh�8�<���V��^u�o�������EcX´@��>���������]�-\Og�]ӻ�Nz�ܿwg����F�>Sղ9�un��H�3�5J�HL��J^�e�g{�`w`'��0WHc�j;c�����='%�4q��G����Zѽ���U�%DW�3f�� �=�J/9�"*@1���q��7����_�ti0(ZN� N�3���23Q�U:]�?x�DONbONu�3J�bD�rǝ�u�B������'�P7���v꠪�a,	Eޱ�V��G8��������B��>���O�S��CO���xj��-!�E��>>>/ٚ��C�+��ZQ��_Pׯ���MNJ�k�bB�Ͻ?��bT�"��u!�18I#�zt������[>V3V�E9����3b�Fg�LԊ{[ ,����nF7�UJ�Z�,YB�g������a��U+?2��tc�>�N}��'�ߝDޚs�e��
�G���Sw�"�ęt�m�m��@
��DD�ޫ¥�/w��X�U(:[�<����Jf�d���[�c{�oJ�_�!o�$�M0n�����gOF��uvֵ]t)((5&�\䅙����/������E��<���p>Ǽ��j�\�V�S�I�_>�x:j`����}�8�G��|S}�Y��~W2R���#��-(���,|�M�Z�|�6�n\��9�eC��'W�4�ś�l_�/��/*P������r<"މ.ej��m���n�R��@P�h�i�H�ň��D�`�rj_n���I��]�F�����̀s����Ø	�������{:��e�{8&Q�H-z��9+��$I�T�>l]�1��S�?��zv AY���y����e%ŋ�Eg;����#E%�I�}�3˔x0���K]���I����?�f�eQ��������k�qX�s\�C�C�%!��_�ō���%�9��~N-ǃ����)�1���H��2��9�p��U�2{m�>+E����PJ���yȳ'�xoSJ�%��;l�Zk�F�Qp��`jf�..�*`��p/� M�.��C��̞�W@<W���g�5�A�i�w��P�jJ4�XCqi����V�b7�8��颚e���z�{2������>K4�+��� S u��p���*�Y�Zm9�њ9�8"�I[���O��s^�sw��3�W ��9a�8Q9��P�<S2v��p��g�o�����n _��-:6�:�;pR� uh'���~�Q_ۇ�q�5<��Y�A]枈-�
���mSj9���w�g:��K1�|h�qNj�^f���n�|b`�=4V�K��TRb/?�e���	2]�N��Ǎ��B�����g,���X=��C:���@_��U:�/Py$[���,V�{]��h�S�R��3��j��{��t��B�{�.��|�Y�G�F{�b�
�2)�I�tş�,���JďL4"��qnM�"!}H�x�UMR\�q{���[5�mt��r,�P&�g}L�-(����������怜�[zY�VR�u.�7o޺��H�=� �ǟg��!P�k=���&��<�8Wv����7϶�����*���P�wA��R���5�&L��y�m�u�W�R�������%�2�kmH��� 28Ś�n���gZJ���+h�;$��G�ҪM2 �+���7w��h�ժ��	���+=|3��7`����ԫ;�:��P��?^�,/���osܦ�4��������=�	�T�T����O�(�RK� ��sX}!׭_Fx.�[ǫ(��.���pB3���S��%��6+���{O������S�q#�jV?�RS�4m5�����;^SƤ$^�߬�O�}����k��e�5��%����K���/��	RsR�[}�#���L��Ig_�w��So�'d�}HSx��)wj��y@*C͖�\of�m�� ����l�޾ٔ��7���Ϟ����i�ĂK�Exqk����Jf]�n��o�frW���3��iϴ�Z:6`��h�u��� ��� y��)��P�ż���{�*k�U[Y�����QRTȃ��U�z�~�7�������?��m�r]S��a��{Q]��~��^8�s�k�A	}{���{�M�H����A���Ky��o���-��05�(+���{��X��t��؈��������I�Z�y����V�Ե��
�J�Y�2�K ����Y6�2��*Qc�V;F����Ogg�#i�i�%�y�!�'���k��i��؂�W�:V����
����ŷg]�d���\7_a���J������jP�#�� ~�J
u[\J��7�u���� /`�������I}�3�BS�E�4Ŝ|�C:��6Ud��D��\�'��������kyԹ��7��f+�@��5��*T�z�l;����a꿦平m�Mx0ބ���$�+�3�>vSAJ4�E�O�ֲ~7���?A�k�L�nlf�>��ލ��7�s�&���#�iW)�}sY$D��֑��D���������S��}�֖p|B)r��'��z^"��&����#V������ "�W��x���-S��Y<+�X�rd|=��[it��� l���0����_���o�����M���E�'q��	~��x�YD%����e��z���K�f{;�~~-"=���e�׉���iP�`+d��=={�T�Ӄ�R�lj���/����)�DL�ތC��n�nn��d�'���h��TUG,���2N[�d�^�zp0x���Ag��z���Od�X��m	HW?֯�e{�-�2�+M�WL�V_�����þ���'���8n�����E�6�)�_��{�ʌ�`*��N2�����d:::�e��ޒ��Qw��0SP�^| �����V+��-ˀ�۲������������	{B���w�S���g5�	�����]���DݽV^��X���oz�+-#c]�9*����n�����:��pB��S���r4=�Ij�4L�raM�u]��c)�,�Y������p�����d���9֕K�i���M(ї<�/?ҊX���M��gl˘��L��{�k
�����("2���i]��"�A���/��,Ŝ�D]H�G�:���Y#�vh~2�j&8E�����DX�&úX
����3���^��٩�����CC.����	oo��|�5k���-�I����.|6}���m�B��F���:L���r�#�h���3�a�S^��֡u���<z�B@@���޼y-��2�~
����h�G���"_oҶ?LҿfZ�����Qqq�ccc��X���b_zu
�-������� #l����6_R��&-�ެ��W�^�]�z�UE"	%7y���l���+O�x3 T@���0��h5��`1��z32��{�j���@�$��X�mslI�QQQ7�Y�E�[$���H'�n�{���Z�zK�"ޓ�PN�^4%�������X�՜Zo�*V��<��L�Zm��F���~U���Fg�AU����zZ"��	,����4O':��:PWf�z6��K�=q'=GY�/	�Ж6�aU�Q_#*s�}���ر�*ӿl	Y������E;�㊅�Jބ2fO6p�A�ZD[���ON��y�[�� �-L�(r�&���z8ܭ���ٝ��O��W�U��ok�l|�.�@���jQ�F� ���u�T}�[WM��&55�ēǏo}�T�	�x��l{~q�3ܰ��꺾��L,�(n��wW��M�cR3x�;�Ub �PWS��ឃy~�|�B�����Z���R�#���1p��<:��:s���w7(( x���`�����VA>�i�&`IL+�eї�uc��N�=��M������Wnb�����~(��s�#�i���� �Jn�w�sC+��>�ׄ�zҳ:�%��8�6KT��ي�ZHo༾��8��;������2M�H���)��솅��K2+�1����ŵ�!{g�ߗ�[}Fir>�+D���E��2y!�����/ک�]����A���ޱ/�Ys�6�$Ѭ���*e��	{�ml��Y�����\Fz_Gp/6�׹����f9��>��,���=!�7mc=uF�OZ�A�-���g�V�
�)�ӹS�4s����s��|KD\>�[�v(�4�WcՍW.����ܕ�����&�D*Y*ܸ�JSx��C�.cC�cC��]�%A�Y��Z��T��ϣu^���Y,�L}���{.��1o���AE�
֋(bn56��a��-jwȖ9#������'��� ���Ӳ�w>��a�Z;�d�A�H?d 2$DQ����o\�Zt3-Mn���TM�8Iw�	_��0�)��y%��k�;�%F2(���)@��8������b�*���y�2�*�$��b��	�馨A����ROe
?E!��S�u����a����}}���]M�8��7^�[�G-.�`�c[~�E+AV.���8���u ��M�==��&Vk�	�@�
��HL�b�ם�VM��WL�Ž�}O4����#ۂ�Bst̔ȕ�5��&4Fý"H�H�,D"|_���(�Nݙ�8�O���+��4Q11�{�Y���)D�#��}��3�������Ӯl��-DA�N�t�6w�u�{�=�2^���L�n���Hiu��*�^�o�A5,�b���F�)5e��q�\k�+@ۡ��l�P)�X�"�`��Y
gj�§g�/{�I�|�[	#�Zo�x[T��Wn�]�i�߽zuI�g���%�#��O���v�w}Fm]���!���D���사o;��$��13�[G3��9K��<���8���|���e�^���������0/�ғ�����Hs��m.�N����=���VW�C��O����H�`�z������'� �
p:L��\�s�^V���^Ip1�:?�t�3g��:Eu���F��V�\�gMd�G��5�8[S��v����T�� g����'�db
�ՠDo�h��谅�A��Z?�gv �n����@V�g��<]ɆӹG��m��D� ���.�]�o����|���o[JAh�g�cx֡I
_w8��)�5�Z����л+��Ar2�#�ց��@�e(�hV*#ռ���B�O��U�ko����|uu�P{��^���/��v$�O����y"�9�1!�VZ���o���c����A胂���2D [xFK�ӂ����j����-C4��ෆ��/����˽y�_��i�0�7�Ia����'���Ӝ�|ш�)�Н���N��)	j^*~l��r�H�Њ�d�����^�W��ŶTT̳�x�
Q�0�-�"���]����#�jV�gn�����vh
�%��V�9!b������EO�D� �	L�=��]tӫP��{��hFĻ�ǅ�)��Y�/'/�&��]���FI����	�KGi0񷘎-.߬��� X��l��M�����;��#���uq�QHG�������Ӧ��F����ER�S��1�� G��Y��Ԙ�ht���ΎPt�Fz�F��&ѺF;\�:u�!Kj�# �PL9b&���#�tO�M���0�AZ�K޽����$<o�R�HÈ��\��e�C����EH`��ю�$���-ے�T CS��6�PS�RJ,i"�#�8_i����q�~_7T*��4gnM�z�����V�6\DDD'���ђ�*C�3�:$�j �'��P������Z~����cd��~F�[o�=mߣ�έ�m�4͓3LN2N��u1��%��NǵAu��1����hO�q��c���n��aX��D���J�M�JC!*ERd'��-�X��=�ІPI��l� )	ٳ�X��Y��X��3ʌ����q���������j���؏�}�g�*�~�?������S����xA�!��Kƚ��[ikA^� �L6	�v�K�c{D�qT��J+��WTT�̺��޻��
C��7�3yM6g8�:W�<Tc	��6��z^c��?F����8�*̌k#��s������V���v(i�wt�x�!��0���h��.�lwc<N�~��!�/ܳ�{m�J,���v�y�'R����	�����u$��FgT)<�H��m���N��^�q��GC��92�������G����4��!� ��>����D:j��Q�އ_�~�O�FZ��@��+t���#M�Maۇ��d��{�3��Z���:<'�f�7� �t�J7�\���ի��fM�!-�6��K��'c�׾/"��y.�p��"�����!g�GJd=�j���r��X������|����_#VA299�nU_��2�����Y�����9��,�����[_w���F�ZoHN�z�2����_��ڰ���?C�@b[vo�7������x�������/����)���*�Z <is�Z�tn�k�U�Jo آ̈}�/9;7)���u3��̽�R��灺Ğw��G�WJ��t0U���v��v�L�}H�u��S�Zp�i��i9b7.��hn��=��?;5��}�7UL�����i�5�$�)܅��%����\\��Î����ʊ�\�^���}غ�9խ�Z|c��̔���}�L�ż�Kh<�m��ȡ���c�G[Qᛑ�-3a�+��< ���ޫW��+�j��>��d�Qhbԑ���.3��8��j�1!�x'
I.�Z�#�4(灌R_�`i�K��M�*�Rr��7�5��Zg��[v��Z{�l���Έ�����W����U<�k���-kۭJ�\c�ꪳVP����m3����*�Ac/��
ha���8���Ӎ(T5�(����#��K>�c�r�C�R}�aS�Q��S�>$������d�a��\C 9y�(e�T���L�0��
���W���:�1%%��l;=&$4� ��� �ὧ�WT��2�cG��	�pt���{Y�؛k}��FY�\�B�1"�X����S+���M�3w�z��S[l���w���e}*�rCºL�#�uu���6����<֝�cظ�j�~J��تl�����=ia='�)U_N��<�Uj1�[�;��g�Y��Z����:�{ɷ޽lx�#�:��������0#��;������мB��W�s.F�;r
��#_6�WdY4d���jd�{��-ֺu�Bi�|0ҷ�X�N|*21D��<~'����m666��5	�0]]]�Y�˓�6#�AO�s��B��@�S�|}M1@}�[����qZ` �U�d���q����2���$�P.'G��34�Š���u3zjF\��i�s����X_ϖ�uZ4������$�	}y�w�$^���>��L�Ѽ:����[������ʶo��������V�@.�{��~J��v�~X�}�tH̺~��UF%�Kݵ��Ͷm/���z�U�u����&)����¢ՙ��<|�F̤�m�	(�1g�.��퉭��::jA�ܜ��(����P+�����l�H��+A��P`Ss7�s���k�����O�ݡ4m�"3�m���{C�t�v�o%Ohܐ�ɨ�\����3�q�:��� ǇҠ��y��C��Ғ1�����%�7��aT0;e#��}<�ۘ���02F�]�7.cVT�A�E*��]�����?O�������L"�̇����%b��[� -�ɘۦ>�p	2h5���{<9�>s,-��`7��9,\�xn�8M8������{Ƨ�b3��1��1��=�L�������7ڈ�Yc��]��N�ɱͮ��c�u#��bx<�lӟ�4�`Z��|�(m��%���ˊ��2��Ȼ3�v� ��jHy�Z=x�y�]Z��Ұk�
�ނ���&�G���ik�Y��Ӯ�r��Щ��/���L�F�]J�Oن�l��A���A�/��d��eDF�<�!2�^�q�c��7��&k�oνC��	��왙�BnBR����p�����j�+���k�9�(A$_�q.˾=�*�9C�uh�l����SN2N����*� 1fC�����L;R�&��P�]�i&}oB��I�G
������K����b�[IB�ΪB�~i��Y��82W���2G��h�Rk����G�і���\)���92U��OR:%bn?x��زu;�b*!����C	�=[�3�!$��G����$oŎ$�~�h��
����	�Ȏ����b�:ߊ��s%߅��v�wd8T�ܷ�,�����|��T3 1Ȥ
�PP:C��O��ʝ&~���D�"J�w�`$U\�2�����96����)�� ����)��+���("9i����Ȕb�����/�(�W��t�I��Mqp�ȈOM�4���>>3NK�ٮz��(�.Q�������a�i��W�t7[�F@[n���P&�⣑G9ω�&c��W����&y��zJr�58d����3$9��[��؝��o�؍�'��GQ�c�����k~��ݿ'%^��G����:SI/� 򤓳�(�>�M݅����9͏�>\ �h��T�p'�1�݄xk/��e����v��,:�l  ��O�\����tv�F���$����<
�sss�;�r@�O�Ǿ���?�*�q����8����bO;��zԞUO���'ۮ�n�t���7�ό����-@��JٞhL��+@��@�?���[ރ���Au�+$s!�3���A���T�r��p�}�@�n,�����A�Z�3�s8w�˳��Þg��u�JH?�$��F>���8 ������T�K_tMp[�{�z��L*p�xi�X������ފI\�X��������4�9?	}y��>h��xiv6�a��i���&�*K\ZA�믶��yӼ4�p4����;�3��f���5�V���#_��zN��Ξ��j�6�V��u��u$zmd/������s���>5�x埽�ȸym���/3�L���	9�Q8��Qڥ�FV�:|Sj	�o	RP�gZ�#'�+ޞo���Ģ�Xj�ԅ��o�?0\9�	GGir�q# sSiswMf��N���u�x�'�3lE��=��(&&�����f�� f�0M�[F��O܀D�� �m��S�Ȭ��K�K���;b��	b3��:�%d�����τ��X�*��P��vA[;^�6�6W?����^��4'��`�,�*��.�Ys��P�Z�{��図�MZp	��Y�<��(���ҍ��nx�t�53�w-�w� �)�v)vhm��.��O/�=?������<4K��������$L���w��q��Y(s�Rs�!ς��u�<8��H�����v�!K;��2�>��+xH�z�T���RG ßkk���!7 TyQe&{��'�V^0͆�:���r����.��3�b��K��"��n`��6���᭘y?2�S�,�잏�}%����1ݚs����(~�v1��Y?_<����Wz�~�z��=J��F�mG�����߶�|�_�9��J��K̶���)=��C}�{��I@0��������Vك���E,�O�Y��v�y'''}ߞ�C�}�87���>KnZs������ޣޛ��ռ/54��j#�ȥl+>v���m᷷���q;��U�X������&���LNVy#}�~9<
G�.�{��[�>D�%Lf?����G�f�Ov��Ef:Y�s�x$
 �c.��H���9Ĵ^Ԅ���ih�&��3͹׬�H���Dv�M���������qNȷZX�m���B7^�6�䀬>�v�V���H��n�`�_��/��O�ӕ�a���R�D�=���s����*�\���9dR���83��(|��VLL�L0�����98f�e{�䳻Ts��[��v��Ң���S+(��g��AWIz�E��6w�<�����2��Y�ǹL���=k5�\�e� ַ|�u�i���[�
M3l	�w�V����*��G����]��D����Hk�5��ob�G�9�GM(rH#PN���D����O:�*Ǐ���x���'�V�����k�á�iߞ��D�<�R{&S_d@��)#$�?ق�x�T��HA`������uϷ%��Z�涀���״�&*ި'�5�����0ؤa[�[�����J�g�we�}���J�;����y{� �w�i�ʍ�>�3������S��wDrӦ-g�.�;�_�:�M��q"e���2}rc��#�e��CW������>S��>���3�S���S�{�Z�h%V��E�Taמ������������u<��=U��RZ�G\^xK]Zs(Z�zu<����*����"�k<uK�,5��w���>< ��������/o��X)9X`O�h�Ki����o�?{����6��
�l�l����Q�Ʈ��XC�k��j�#Nn�0*��`�v3l��/�"�["����u'�F2��v�O���Sh^�0$G��>�p �|���=yCo܆�����氝������}N��[26Ykf[J����� F_����s�}c 4u#��?�G>��C$���_m�w���t�VK�uz���@���0�#i��l늛ɇ�0��?h4)_͌M�g�f��]Φm۶��>K�y��-v��(�Z��z#�-����pg��]V`EIf��p�1�j���QB��s+LwY7�l�u�W��{J"�Tȉ����ꟄQg���ض��Z��xv����^��mKK�D�� �nn�����6�J�S�x�Ίt4�ewM��A�(w+�q/ܶ����hB���Z�Nrzū�~3�ES��b�(�ݽ��=M$21a/pd���H�,,'�=]�m�r�wP׀��ɭ+T+�����Zw��c�]ùB��/��R���˙��sr���]���Qq�N(.�.iﮞO�L�Ć�
���q�{*7b������Cw�4q��zQ�[�#^��9���4�ar��稨L�yo!�A0;�Ѱ�}��F�j���Euv��ҾO}�d���@-��\�GUJ��+���ju��tސ�4kK8r%B�6,�mz�T:��c���:��s�c���)�@7���ˇ�um�"}��G����]���x���z�a|]cCΫ9���O�e_�*���7��e��e)e\:�z�����'&�g.��dL�Ĝ_��Xb�Uaw��]=�3oBZd�=��_i��葧�V�=���i+ L�z[*[��Ťq/�bK��L[Ǖ�'�B�l�Wb�n/�Z�s&�\�qZiw����Cϖ��Im�+�׬��Q��-d�hR�z^i99�܎�V�f맀���(˃���� ���	=��6�C�~��ɕ���o�
x�z���πUT<�k������pj�?c�ZdY�S��7�CEzsUg����5_����G����h�7���T�nk�R���?�4�$$$v��z�
���$펣�򷪩����0�/�-6J럝���+	��F���n�$���8e$��S#h��^��k�Ͼ�S�"ɮ���٩C���y�<���>c���7���|,�W�����+/�!1�Uߖ�%	Aw6O���]N\���JJ���K}��=�0������\LXBb�u���腓��a��Zl0��#>,�!`2U��῏6ښ��J(�D@ԁ>Ź�w�����4�6Wc��ל���{�{��K��l������'##��d��hT��v/l����֊.�Z���!���oݖc�m}q�����/���T���0=��fn�GLl����G
�X���6j��$O������^P�����@
��{ai�Ӳ���f�*o�;�E-��{q6<2����$�R��3CV��R��V���ޱ���f������3Gc���b�{7��P�%%%�[�^��+��R���� �����ߖ�C}�
o�p���L4����%|L�wҎ���k&j�
��֥�Vy��H��F��	디�t��@$Zoo����ν�P-9n4�l��&�+�1����Z1&$/:�+2Ya�N��z0�|�O�� �4Η��fĆ޸q$t9��.�'2��)}�3\�T糄�m����2���켦�`fp�&8�F�`�T/z��Pj%�]�m����g�%�VŻ.�1[�L|�릐�1��ϫE�L�ȭ5����A�: z{�`�aվ�dh}���	k%����|-H�d��s(	�x�>�#}Ak��ڃ���C�pB�\��ǿ�MmFF8r4�CMe��K�}_�K�i�U�ׅ3�L2��
�[��ǟ;@^�A+��x�;�OE/�r�Y�	�Mqc�yJ#nF�V��	5፝�q���nP^����B:��lFRC���*�w�]﮻����v���®U!|e:�T���5f{<#�x?�ظ�k�����sww�Wq�[�ѳ]2(�T[>��LZc�q�ZFsP=��p��`kH3��m�m�Ov��#>����/��`S���t�cԫ�*��i/�)))�M#�K��[9*ja��U:��4d~�eR{QK6:�XV4MV�˃>��W�6�;�@��]�������f+r���3���g���l �����g-�^�Y��d,��h�����@H��Z�D����1�H��Km�S%G��0����T]l/���{��M���.�x��� �Od+kUVT�$�)�O���hKx���l_3o�ծ�"���j���[�]�v���	��������X�ۃ��X�h��{p�b�Aa���������A�s�p>��?�/ŜTn�	;��V2Z=Wf ������&�455�𷆉���VnԢ�П�����Ǽj�򥏏;�T��@Q��&�ꊸb�q�@����[&j��6�"�[��4��=���X�zG��>g{y�x�Зh��|�K|�o��'P/{)|�����1����A�-�~���dꇺ楴����h�oJ>��L'(v�ϑ����ϕBҫ�>��O���pjz}9�Ou���3���d-W���s������������[榦h佫����3�f�g�Uw�̰��a�`�)��i`]m,f�_�PU�?�7ۊ�jn����O{A0�t.�.oz������h���_��3=>���"�ʄ}�Y<�C��:[���,�ƽ=�u��WT�����cgg������1v���O��N�*��\QYك�׶	����ٱL}�@�:�ߵ�j�ѡ<��U�'�bX�5�$��&?�L�Լ�*�A����_`Qyy�zi����]1���+�P:r#��g܂��v��1�k<p�*T��k������C�[(�lAig�TRt�u�#h�%�K�Kk%�묐����hC�/�λ�V*����] �"�����f� �������J���üw>�9�8�x�7�/��|9<�
A���?�y{ T����>;�����^Nb�3�qH���A�XgF�B%���wbg+f�����?��tK�ƞ7w���jIy�[��vrsyv��U����uǌ=�!������I�8�6��O�U�6h��rkZ���	�c���cB����dM����ܹ�	 �Y���ޔ�oZ�P4��N ��NN�և���B���������A��Wխ�1�7�B�&��lB����&�L+E�zA�ׂ���M��2%�[��<AN>��E
i�^�ۉ�9t�B�E�Qdٕ����h��%�R�i���v�L}�0'RO��(��!�P��[U��� �G��S��_bvP�����4�5�hdbvi���Nhyt��Px��ir�e��T��+y@V���ӝ���#N>�yMg����ʕe�٢�ۭn<�מ����н'�=�Ѱp�Ҋ7�J�N�g$?����J!��yy�6��L U~�,�J.�|S�zdd$����QQ���kNy/@#L̗n��3�h��WV�]��O�Gw���@Ko���IW�$�?��'X@	S���6��|ҹ[����.��1�Qu��Z���=9�y���G#�B�R��f��v]X����6�o�}b���3yLt�f��z���ҍ��T��������G�}A���U"h�W�J���Аe�����5�F弁�~�=�5�8;��/xA�Lڳ�g�-��>c�Ƀ��Cb���b{�=�7��V�У�׹8��)������)_k���:��+����n�(��L�ι��>��XzKv�� ۘ��!�b?H.����G"j��L�܌���O��m��uR�l������j���Ɖ�۷-�v���ˮ]#�B�ڢ���Wȇf��eŅr*�؅�a�D�[�lg;%ona�?R}�}r�_�lܛˍ�
����lK���K�K�[�y��  ���u�Nk��-3c�o���N���e��' �Z] ��_ܼ>ѝ���M$�Eb���j����h�Q.=��ܤp?hN����M
tk��_Kka?�o����M}���2*�������9���T��Ƭ��b��tR�$�*��2����U�' �`�D^�~%Yp�޿�qv��f.%��DvJ鰕�����4/�@=m#3*����|��w��Fy���^٦�
��V�����YТ���O�U�V���P��|Z�`���d	l렱`�m̉X�����7��Q����A'��h�)k�����2F�O�+/�.�7�Ko�zv,�DN��\rȀ1s`rD1��:��LDQ�R����tҵX:)��t"*V��_�>xb���h�6y/@C-l��>�F���'�֗/oG�JR�)��4��D�444�-�Ux�S���/�,��M�!����GR��̝��^���ɠ9��e+[��[5Q�Px��
��ʴ�$;H�jz):]�Wx^U��=�5C˗@���;i�-��.�q�'nyS�^��1/r�b��)5#d���U8C,��i����� ꩏�{��e k��pc�./�j�N�����%9(�6[<��
9r�/n</���[B̆ٶ�]������^�#;�?��YA�t �d�R�V�b_{D~u��[O�����'��]ŋɻ��ן			h��5N�ʔ�;��#3�m���u]l�T~ؽ���dE�ɧ�CM�&��֙���c�A�
]�od�ة��������;�pB��bq���]ba2U�2u����379<�9�����K��|�E���6g1!�@H�MYW� W��?���䞎TUS�)l�[0�Rnze���F�������j*L���q��j0"Q�g�H���>���)�E����ǱJ�R0Н��A��'�9��!��Q�O^�ѯ$F�o�<ğ���Т��Z�}�Μ�P�g ~zr���f�m"���W�}�������]9<���(�}���xm��C��3�Pd=�}ꓯٿ�u�r�_��⎜��)�������z� h�>ߤd�?��P�s�[e+6��,5_�S�5�$�v�B1�<����Hܕ�����F�XR���wyk�s^ז�f�k�h�ly���5Tl������m�k����Di�L�����=�����=��g�U9�w׻%��D��yV��[�ALn�-��t��=-�3H�`�u)m���j��64ҧ�= ɖ���J�����2�p'!�q;���>�^6�9Q?ŵ�#���ѓ�-dW@����i8�͈/�gђۖ6v>���>�V�|�YB��?���{�[La�?�ح7~���1i4'�?F3-��pi2��Xw
����v��r[n2t����3�)������P/x��zN�ȃL"�r��2f��f��Ta-rX��9F���n~皑������,��	���]*u��^��ڽ��&A�����������>U�ne����d�Z*�!݁�ꠘ^�<0�Q�@���f��>K�s�6��k�
ɕx��FQ���
���ԡf�a�RTg��T�%E3��/Vl�y�4I] 2�^������}�5�+
��TI�l��~�����Rb�,��p�ؾf��#�~Ʌ��Ùo�
�%��bD�{Lv$"�sk���H�iɝ��T���OQ_�$'q?�bR�Z�:����ڵk`%�O���C_�t�|���A�on"ln]�̐���土� OؤώFY9��hN7��y��z1��3�ފv���L�2����=y�g���ݓ���U]ö1V <=�ȿ�w�"###���A:�.�xi~n<Q1Tӳ��!��@z@
���Tc�����ƒOǇ�V��
fQ��A�V�<r�Ϻ��E?_R��:&h$`�^n���לām��%�$�ccc��g�c�њk|��n��5̱�,2Ѩ#��$$$�<*�|�H�l��[Ю�ޕ%|������m��1�ݪ03�Y��?�@l�9�z.K؁�p+��+����4�8H+/�V�0�͝m�&W	�4tS�:�b�<I�)�
G�����B}|�#����P=��s�Ö��|�err�56A/����x��'7~�K�}/ =��:.�׭� �;���P��$���������K�y��?ޏ �U@&s��U�������v	���#X:ț�h�������e�E� c!��t�0���)�^��TyZ")+lWZ��pէЭnU)v}��A*����:�Þ�����k!��l���� #��9��㏎w1�j��;#ܾfĬAJ�2��z]7 ��`��)t��.;,v���Wy"3�4������c3��n5�����N?ƴ�����S�:�ȗNt/��jMLL�s�(2�!���;�2�f�݅j�� 9�K:�d�f4x=�65�X�n2U;�>zh�U�G���S�z����4���C��J�V6+,�� �aA#g-HZiQ��[k.�K9m�л�t���R���6ۃ斖���0:� _fڶd�V���D肐�鎠��Ki��f��n�nod�i`h`���[T�	q�icO���h�󚴗�v�d���P�|9Q�On"��j}A�ò�zF{��	F�8�?=*�3�zf���ߙ����"f����V�\��!3�8�Vg��	��sf�$�h�'ɽ�Pu�̡�f�X]#���s�Ua�{r�&��U�R~�ICquN�!eZss3���-�cMf��d��Њ<E<Ri�%���d�L�������uk�@�ɞ��]c�(/w.�sa�PlYZD K��YK�j�A�����8�drG���]s�9�2�}ޕ�H��3�`�q�HJ�XJ[r�c5�Ҳׯ� �BN&�h7�kefg�Ǯp�:A�.���WS�>E�{��rn��4[�Fא��W�2c�/�c��N	E�'��{C����#GX�9���rmwrƗû��v�u�\�Fz�� ��[	|��g?#�����e�����?ز�F��pPϾ�G"�V[Qq
y�&,��߅<���Ӻ*4�=; P�ZMlK]�]�=�H>���x�IK;E���E\�|��W�k�Vŷ��.�D��D�B4@�T$#E�(B�%��W&V�ʋ�aޘj�n�6y��E`��?f��S
>��R����l+�|qEz`��la�T+3�hp��=Ə*-�[6�<)���bgh�b��v��=�9����5t*9�gA�*���/e��5bv@ü��E�����^�VL)����{���b�g����66��(AO�*��&�O�~d�"�O��s�z#����LA�����:U_Cb��%J��ͺu�Q�D�)W�h�:U��"L�)��V��n�K/�6`�n�z'�c����.�w�)Ni���fF�����w�9����Rf\)S?T�Z� �鱪��{r6"�#�B��8�VK�"���Q��ҡqE����	d�FCͯfv�U|F��v���w�DD8;C�R���*"#<�6����K��2�%�IH �3� `�C��y�RJk^�Z��������,���ck`��e� ����'�s�3#�ba1n�{��d���B���a��[=�eU4�����F������V�^AQ��RVx���Ek�qXH��P���K�P����R��5��n��	C[���0�(���C�,.V�)�w��t$��Y(1�L�� �,�Ki�-,���\��TQEBv��.^�����64�5Q�2��ܽ�{��뗼lz����pӜ%��Z9;�����q]B%�a�;�g�ڵk�A����*��z�_ `�[���l<^��5�=~�b��zB�P4ˮu=t�Zi�X��E���i#�}�>o��`�2�ŖS�m�d ;n����dd�AS��3|��=U ��
k<'ɣn�����m/@#�{�&U�v���۪��fԷ���1.�u����\~��cQ�RO���"*=��f��eU��ٶ����ybb#4��6U��G�#��ѕ�U���^ڕq���T�I\Y�;l�X?F�qm�P�ɏ̵ٗζӠ_AAA4T���A�K�[d�z˼M$�&i�s���J���o4�z����n�gEp�2L���(�D�ċW�f�]W<@�y�s�N������{Aydΐ���5�ik0�)����A���h���̯⬙�Ʌ������v�5�"�r׃�M�K1���MM ��
��n.��˴w����\�EVn+.e�=�gLCK���[Y�d�E<�~A�CZ����v����os$��Sq�����^��h�����)������,��ĺ[V����~d��������m��_��8���R�ˮ��� JϾ:�j����b��E���U�L�@���[�+�S�R)���6�Z���S�)���R����+�6��e��T!�.U���G���E���W@�E��i+���o�Sf�n�\k��}\�j�A���W�D?ʱ ����nX�?D��� ��-����)�<x��D�
n��oa����$nB���"�'�? ���-t���]֐?�2����V��C�_a�~�l��>���r�sf}��|��m�)�9u.����*ր�����I>>��MwH����у"���ʾ�щ�Ӡdy�)�/Kyx��c?r�U�u>u%�{�Ү0EQ�y���W 6�y�( ����W�B��q���7���f(����Xf��
'r��M�3Ya�o�@��w�@J�2J��aZؖ�V��64��Ҷ��� s]{�+{���W+N��bW�8Z?�3�������y�㷫�Om��Gmu�}��("��s� �c�x�[�mv]k����I��՜j� �����*r���?P�����C��4��^	d��W��mt��Q�E�#_af,��`g<o��'�_	�F�+�՞w���{��d�>?�m��Ԓ��X�~�����554R���^@�ɼ���Y)UL-�3W�>��MrJSS27�2��E������R�z<1��U���Z�۪��z�ҥn��6�̳�!�{U��L��F[��t�ڲͶ���4U �����p�{��A�*׷ɱ���Dy:�� ����9!��B�Ѐ��?nV�ƃ�v�#��i=^�
uۮɨ����J?�:�E�7Z9�ЬjܥK[�������L�\̑3"�X1U�qͯ:�U�V�s;����{��=��x����3�>��k7���uĬƇg��A��o~��p"&�9[fc��B�x��N�C��R���b���B�e�1��db?ڋ�������PR^�w0����ylk9��y���_j��K�>��7�B���>��� k�8��Ir�Z�h�[^4B'Ś��p ��e�/�H:���ޏ�}�l�"66��/�-�q��.W+�����?҂�ȏ��^:��Xt��ƶ�a�0񗗬l���
d:��&��ݻ�/��_P�q�9(�%��#��Rښ?j��mD�}�����5mVi�M���㘐��*��K�)f��/��Q�B��-����3��qu��`����@�G�U��i���c斢'�__�%�C-)�qX�qT�����V�]u\��POe>A��_��nrҶܔ���VT�����c�=9J��>3woϼ훕h:�k*-e���+������s�V��P$��/R� �8-M���ǴZS��}�_��!$��w,�al�w��&�E�n�a�L��6B����s~Y���&S?$,LL�=k���٭��²�4�_UQQ��i�z�����<�=��]��Y?��ø�?�O�뱔>��1,A!���#�����+�]]]!�e�X^���6�R����L��"B��	��>p�����B j� �6�A�jv����ה�PΐNB���4$Zh�ͱ�;�jb����}��Xf4�\�g�]�h�RڽyW�����b�cŢ�J^��b�4)Oe���BBJ>}�4R�stt�$�p�3��$������¢���y��9HX����[>���63�4���&�?c�����v8/d�Hv�͢I�bU��o�B����`fF�#Fz�� �C�V�,ha㼩9H�6#�y�/>��bw����B��������N�1+�N���������2�G�M$�.���i?C$)_l,/>� s�#���_N��:~�{6�38�͡���L��0���*"lD�?G�����)=i^�IN�JU���x���Kո+Wv�Y�s�f���+w�A�f5�'���W<6��9~��jm��
n�)�H�{>$=І�1��@���a�7�2p��C�o,�ud=c�[E�K�\q��B��FGWb��^�Ĕ��h�"��y�Dh�1��4�c�/e�)[%�5�+"�z��/�3t��ޗ�z��Ϩ�_�]��"�b7*�/�g;�2ڌ�ȟ����V�$�?F||�{�"�oa��y�+�r�yA��:k.?v`*�-c������Czۿ>�02& ��a9��6C�:ɥ�-��m��l���#��3��7��$�#�A[�8	���j�yΌys�x	�����[T[��;N�&Ă�q^^
�����+/Z�`'|�/���yO���2�uL�z2>��+N҉c��FX�Zr3Џ��k�xY��1�[g�)�Owh�r�Chh u������|�_�B�
=��7/^��Կ�����5[qji�<�����<3';4�!ζ;��5����l�ݒ�=h��k�o@_',|��]�v�M��ŮSЂ�B�R�A�]��D��)�'�Ȭ�IC��Tvc�]� �h�F�Y �(���t�O��ѻ9�;�!�]�:���p�v-V��1�v�nElY�̞�_��A�Y|�A���"����I������]�b�=���"k��
(��7�`�z&�x������A����ˋ�������
�wv1=.n=���{A�)f.{��؎�p�C�ńz�Mp�lǿh;�(�
�,�bV��x�C�����ȜY��̼6��|Q�N,��Zq�"aq�'[���y7�=���� ��C�p��M5������a��W�V(t���b�	���e�S$���-�_ͣ0񄿵����ҁ�Y}h�ө�=%���Й*�W+3��ļص�����y6g�&�֭�8de�� ��.�T/�cy��&[���+X�!�Ӵ�e!�
3�%��,�<����E9�2�qe�I�eAN���A�b@z��a�qA_t�̫� WO�����tL�Y���m�\,[n+vݾ���*v��,���Mj,d�W��`�)2x�&����f2��� ��r.d&�Yt��Tw�������H
�KZN9������t�׋D�=�d�������9ʾ,d��2Cqm�E�ca����?G9�E�f^����,J:#P�j*�g��k�-��f�%,�|b�A��� ����	F�߯Hdł&�Z�Nj���D�m|:��'�5�J7�#��ψ�=�˭9��Hg-�ޛ�$�	U^}h�&���^Ǥp!䵈��;��J-B�E|\�"AU��R-l�#/9����_�\�G�0����jzz�Úy����Wr����r��-{lH�d*a]�k�&���>sC����
��4ˆ]�����9���7k�V�� �o{�Qg����F?,��e2,�f�}���,{$�ζ��{C�;��P^�];@3�����,����F��Z�l(�Bd�p��;���-@6���UL���-���;�C\�u{e�Q{�]G9b�g����Ng�-����1�s�{ D�5c��G�V��,1���oZ���2�	\�l7S%��}/��k��QE�.׳����kX�I
��Z9�?g���%[���w"�c���p��H��
��	�L��D�Lβ��L%�����7\G�ä���a�'���JX(
#�;����(l�L_.2����9�He̋�AK�U�?62M1�.*17t��g�HK�2}���鼎�D�"��#a�DL-�\_F���G���BtLl�&������"�/}c==@w��{SSii��ϟ?�gg0����T���#�b�!�O��%��c���u�OHp������_[�s濎�+3�u�ԁ�3�u�|����.�K�/����K�/����K�/����K�/���O"�؜i.���7m��W%;+޵�ؾ�����K��_#�_�	�%���_�	�%���_�	�%���_��oߔ��^�����K�/����lo^��#�^P��!�@���H���/l>jB�%n�����X�Lŉ�*�?�,Y��[���������}tOt�H!?��5��%���i&�}��c�Y�s;�u��b�l��r[�g�����ӏ�|8q��z�ի��9±�sS��D��Z�Q��b_r)s��ت�on=���r���e��#�.ee���E,�W�*��rVY�n\��|Y���c��Gi�/ɿ$��N�OY���p;w=�7��7�EݞP8������YZZ~��}�����W�P���X6gX̥��{��_�I�%�� �EOW�3��S�RZ�v��ֵ�Y���R=�P(zl��ܴͣ���`��	��-6i3t�C���	�U˙>I�5��TTTx~�L��~�,����P��{���&,Oz��5E�$Gxs�v)�*�����#�����$���G�,]��i���_=k�����cy���Z2���ˀ{��>���d�f���.b�|��m�С?6~���NؗUD`y&���r$i����ٻ���0q[=v�c��_�	gw�A��g�,� vJDh���=���b��m���A(JN���t��
M#�yR���p?��������E�Mp?�?V���Ս�%�8k�2�Բ���T�{��/�[4-�$�J�M��5��-t8��Дm��b��r�/��7�Ȧ�o�OG��C;rrZAP�U�����W��P����c�lj(�������?zO=��t�j���
g�]�V��^h����M����>Y�����0NR���yA�yCYk8�N>+&��b�/�)Ύ����F��G�Or:�T����D�#�Ί2�T�~�c^<K(��f��k�CY��ۙ�t���?6/z�A�N�ӑC��q���E����ͬ]t�%'�T��K�U��D�B/���pߗh����"�"��5)�-�I�<8�v�j��.��Ҽ]���OQ�S��('X��q�ys����pR��oXm���8���J�Z��:�A*=�*]�V۴�"��E7S�S��ݠ�ɏ�p�y�%��1����o���g�ٝ����U�y��d����9�0�]��%������t��r�}}� ��[,����.}�>3=9&��{0��6?���&8���;bXe��lj�\J�c%ݽ�J]�#�����m��b��e��`///w�2î�$	��|$JRJ�tr�y�׮-_��aۑ��#���#��R��yw�l���u�������	���	���G���>�6����n&+����?fX'�@��~'�7';�EV��Y��[�����GHE��fO4}Q]J�Q�;�fMJuR�S�k��D����������+}�j�r��fh]�yX�}&x����S\���}�o�Yu|o��U�r��V%����m#�]�C�G��{g����E��4���[m��SHwYe���"����?��L�-�E_���sV�^��\)��$I;я|ʯ(Z�y^�y�#ފ�p��bד�9�,��P���E�����a��x��Jv��q�E�f����p�rʩ0Q�Ul(�Nm`1�������U<��&9�e';4x����҇K��fr�g}��^3T3'i�%�Ƒ�r���MŮ�:4�����6��rJ��?�5��@f=���zFF����M朤j,����������Yu�bjY�<�6}?=:�/�nݠ2�M_����L% 3����X�_o�2������#Ĕ�ԏ��5�1!���N�yi���A�癟S.K1�V�~���8�����N���[�!13�(o�p�n��ЄEЧ[l���s�jX�Sq[���E���!"\��{��U=����>���sq��C��ܒ�
�sd{oa��������&��ǯ響�K�,���\~���ci�����s��r�g����D�q�L?��:?C��꫔�tp��PU����g���)��(����ut�����y_�E�cԞ�ư�q���U�j��a���Tc�N�����qe�=u�:�.�c-���߮rw%!�+��������ͬr�qw�\��? �{E��̔K�_�e��	�5c䅒���?��	4�_�?�+
e)�!��";�%B�"��I�ƒ])�P�]��lY"	YJƮ�e���wg������?��;���~~9���������}����˹%���TJ�Ԁ*�7G�r�\�N�y���Th�8p�S;�]���߈�H[M�zQ�2��*��`|O胚�[h&�R�n�T�9�f�Ǽ59P3���{N@�m)��>M5j���j��������ʍ�oXX�aнΚ�Ʌ�rBC� vnr�B�(Q�96��7�	���A��^l3�C��"m}�\�Jֶ����Թ�P�?p�R0��Jc߶)�����r�*)K��N�FT���˗AD�S�\��FY��������f9�C���i :6�댧��Y�����a�s�s��q���*���V[+Q��ӯ� �"B��K ��iFVy�Z��ۣ���9�W��S�4�W��=`��Ete��5�A����� V�A�4�LdyU^j�����DUy}E��|�y	ç����Wq|�Ty�����S�` �~/�a��(��ǩ�J09�1��B���6�WXU�c�2�^^E�F
\c\U�@2���t�`ek{���I�c6���<ԉ�݋�{�Ʌ�{>C�G������ ����6'��f'�:��Z�6S��~\��T��o�	�*s�Ǧ����J�㍴@��_�����xsE��-��&C�ԣL��+1T�2���3��h�.��m+�ċkq��f�|!y�D��[��p�k�c-g���ʘ�@�e�ktR�d�e�����ӧ)�]�Z�v@>Ń���� ��0�Q�j�B�Jɛ�q6-k��YB轚d��i���r}��J� ���|1r�u<q�7�0��� i�cةAS�bWk;JA�i�<v������f�٬�E�>�c�QQ��۵�8%�ض𽋪O�!�Bwv��ϑ�E	OSc��z�u<���q�6W{��e)�zP�vc�D" Q�c<Q�eO	'1��x���mAx[z�n|�|Ϻ1M�U\�a��A��E�SԈ����`8�W��۹ �B8�[���m೟��:�ǡ�ܲu����8�*p��[�d�-��W��@ʧ�ĳ�� �ߙw@�G��Fi�-a�*�����^v��E//����.���@B'Ū��"��,Ÿ�޷� | �A*�����Y;������}���x;H���K� ˴K�:}��]]c/�@�w��p'�7���pY
3�]�w`�d%_��!l�v�WQ���T��+�~1sq�D��4ŉϏ���(`v�p���p_��;y�6#ɛQ̾�������[�êd<gj
�^E�i��hli���/E���
�N�&?�R��󘪝ȫd6σ2P�+;�q2��w�ǳ�����ۭRɨ]['��4��ߟ``0sp8��6"���[��'p� �O�b����_�VK����Ē�ʋ�Q��_{�}�=�0��T�r����_���A�ҿ�ゾQ�r���dA��Z�y#'Z>_�xA>q�W#χ=��!WO��sӞ�'l\d��)ɥ��q?$�^�Y��rvш I��
Pd\u��)��_���T���-	))[�(K��4�N}T#�r�毈�y�:���W����`uڈM%�7Nmی�o�,�XD-W<Cy�����ƒ���HR#�����V�- U�dS��ڄM��ZaF��m��r3
@��:pQ�� �Ym�m���j\aEU�2Z�?ΕǄ���쵻�f�1�s=�5��:��>���.b�57���ܻ|�;~���=�l�	��mD��z��J�~!@)[�K6V6\6�~P)�I@P��+iMH)����5��3�,zm�7�:�f/�j�NX�-��Iȱ�� ��.y2���%��E��l0��p�5�l+f|��.ӧp&]���am���/���^�,n�7�Y���LR�,��0������;),�I��!t�7�Q�9�-�����Ɠ��{Cm��j��l�$V%�-;R��� �E%����[�2��5�0U�i��4�[S�V÷�]]z�?^�48��ɬ�k��!m[���ON�w��l����#-ך�W�8w�f��뭧�$���W1�&�����GA7ϝ����
�s�4}�KgR�b�d���xI�Թ´��1��~�t�)�UKjp�=MAP�t_�����E� %A�jqi?�;U�=�N�&Da�o\�r3�
BMx0�:�M�"��kw=�PjS�*"X�����"e� X)��w��0j��pce"ovc}��`��z�H�������D��TA	O�b�v��	�Mx����8Dx����ׄ�:��4yC3�CJU��(:�	:���R�����%0&" �"?@���pV�k�1᥹�pI[�=��;]G	����:�MMpD�:�"��ܗ�e�)��Q�$����ɇ�S��"<pJ�R� H!��c�,����s��t�{�dv nH�u^KGG��P�ˀZ��nr�qWS|+�)t��N���� a�� 5Wq@P�Э("]�E�nܬ����J���!<���
�	z�E&���+w�TH~tE�u�0r����ՎoP���+|6��{Z�A�zSְېǂN��ѵ�W�<���jb_,��tA-n��I�xԆ��S�Zm�-�;@�����S�{ �$CW}	9�|k�:j�&�n�N�T`��̬�����^;n�z�/r�F��
)564�h�"��A��zp��S��+۸`� .k2��� N�R��ww!(uR�� �	�#�1�;]����C��EU��YY_�Oڐ�����ۦ>,	8�TNg�^���>w���9J�$ ���B�A�9���)P~��.��Q��I� M�h�*Fs���G%�KiL�|��2~��r**-+�~N�]���cH��@�U��u|dd�T�k+XI�"ͥ�|(P2�_ö��9	(􄅅EZ���x�/�lk`F�6�*>�7\��_�rC(h�,�����p4QukN�O���[��i}e���01?��a�v�'&�G�طf�*�>'J�4p���ɫV�ǣ��l5ǥ��d�Ȧ&�~*RE
��DGG����.Z���������l�P�b���ѷ��@J"�ڴ���n���X_��$Y����7�����|cl`�tC�rv�@9j�`@#Oݻ]�XH&D~sԋl4�5�|[ 䓡I��=���U~_��I�:6�[�4aa�ق� �4��J�բ�	���K (^�[��A�����IX]�<�kjx�qdnv��*�,���
F��5PW�������#h�׋�Jj��՗�H�C,��M�&A�o�:����_�u��O�j��=� 4p$(�"��+l7d$$f���Ń����\:�]���Rv�U�Z'�0HZ�'��Wf��7eFڈ�x���/�����bǄ3H$K�l��l��j=[�'z���=ѓv����u���_��u���_��u���_���w�y�$��ՙ���}L��� �/�9t��BΑ2��
��)�n{=�͝-3�Fg�y�?�	�~��3��=y�!��]B�"�S\V)�2��R�˛5�@~�<1zb���Oo싳�X6��X,�K�߫���}vR��:%�6=��4�Y�a��\��~5�<��`'�,ƶ�#�L�97���TO��TR�\������S���-���uӃ5���*�����9e�f��eW���)�{^Fz��ZM��n~r�n�h3"��2hUW��p�/2B�b�ݍ�"�OH�+a���f7�G����CL~�CNU9�����{�AL��Y�ʤ��{z����ک)C�#Ĉ���>>fc�	�'B��@�[��<���0���<�&��Ջ�H1���>��	�q�F�X�����@�8|�Zg�g�Q6�������.r�\��ַ$��Z�ʅ���::#�����7�j�e�V{F6�֮�8x�Kߋ�̚X��Ϋ(��8���[���ה�̦̈��"ߎ�!����of=Wڒ6<��-��A������/ ��F�;Iz��L=^����?��	�mw��/^��X9��)�D��Q�h{/�R�)`��d��k�5�F1��潧�+������]൱-I�=��Q�ξ�s��m�/���[u�un�%��Mڥ�����jQ��r~��Wv���"��������V�Q��s�����__$C�m�/洩���$��L�jQ�`&ڳ��?9���Md�E��U뻉6�W/6�!�o��|g" �&"4�^�'C[%܆�>P4r&s�P��|)��]�&z*�?�� p,I�H��kH��;�N�y���A��H��c7�5��Xvb"�IT/.� ����Q���q����!���#�m���<�N�T/�iń_�!�P��3܉9D�V@H�(&��W��PU^K���Bhŧ���뜰�����Q�;K�s��N��>S�k*\6#�;1,D[�iM�-�)�����[4~���!9����L��F`�*NJT	��PH�Jg�-e��	B��l6#�d�3�/ZT�S�$��-�[;n�O��U%0n��7�F��F�	����L��&�-m�?�
	��G��e�-�u%|% ����	&���e��z���.B��:5x������T��8m�c�a�� �x�Aw�Nf��ss��� ���4~/�>�ᠥ/Ҝ6#C,R��>kì�e�e����F�Jf�A�����?��.��f꿟罐}����5(���<�n\��1���ߜt�(�̐Y���^�tIp�Gs|2��L"	AI�R��_/�l8"��'P�M�����
�R��Pѽ;)�YO.�E����i��qy���'���D\�J%�6�)�א���� 6*<��=��*��هp�f�0���LQ��y@��m؇r�i��M��c6�i�`�mƦI+�oeM�	���?���*��I�b�,m�K�]���	_�v��f���vV�&ܣA��`.��vBK�~�v���?����`�����4+`/+03}`��Χp���WK��4'��0-��EE�?l2�l�%̾6 A��O����qF Ũ�Y�?�Iıqh���B�a��9�n�`{Հ^���j�z�;�Y���J H�b��Mݚ��g�?�=	���t����M߀�B��k����8�����U��w�e�Bڢ~�?�?N:�O#W��|�+7��6q'�_RH����@��񭑡����Ǳ�:��"���Z�e��3~�T���j��IA�VO��R��(�ǈ��aA�}-,�1�y?�eʞ5�0+=�s�#E���Zdq-���>�?�P���9�W� s��N�;b�<=�3[q@�1h<��c�ߡ9♕���Ǐ/=�h�2~��bhq-�* ��f|����o-��P��G\�3.����M�l|+h�%n�0�ZR�V���H��a8E�e�	V�b��j�cDq#+F����.����:�<��@��/�L`U97��7�qс-!Z�����k)�$���-��q�� ���Ȫ���;��8J��s��D�Q�F�G�hN��&h�Ǚ���NĂ`P\�8��t�U f7A�c�J�p:Flu;- �q��]�T.؈�}VTp}A�C�}�ذ9	ZB�#q��o.-�EO	�o-xU?�▢�}({���yz�𝮡�A����nU1h<4�c0�ߠ��吡���9z�K�T�8�����=���8�����9�o9��!�z0C��p��;���b�'C�%JT��0XQ��&�uN��^��:"�n�-]A�h�%�+n�P���2��q} �U	��t�� b����N7������H��}X@���[ú6@^���Q��D�,ۺ���e�-!=��&�Q*��Z�}Qo&aʓ�T�#�[��f���_��1��P���"��xc6jf.i�L���z��S2�V��k`�������4 �l�ڍ�V�_7����RI�3,u���QF��=�
%�Ԯ�`u����F �P�������.��׎!�����m4>+�tRݵ��YY�-�5��0���0Q��x������3CK���z�fP�r��ZF[����)4>�
���)�xD��`Vř�K���N�_�C��R줎b�XWT����x$��å�0^#�gk;�S第�˞,���YYRԴE5�=�`��*��,w�Ӯ���S����8LP��sM2�{�9%����4Pe
R,���^�XB�ʍ�K�A���	�(uR���hd��WX礋�d���>[ߡK:��
T���Aa�	8C����)K�8CdA�ݰۙ�[I��Q ���� :�wD/�B�
��D���!Ga{"��F��7(��������������s�t���f2���.?(�Q�H�b�EѸ�)��8��M�
u{b ".X��?:��?�6���!�"y(Ei2tD��^{u��F���dC2�c`#��������]nr�A�eG�%��s�T���kŨ�1x��[$v/���[F
��=���q��f
}W��a�{h�l	BK�~V�>��Fb`�I�':R�0@���ԉ�ݖAH'A ��"��R��v�r6�s)����ʔk�0�G�V�Ƅ1���:�{�+є:]����7�yr�;��A �-ub�ODO~s�J���Zt�{���\����3n����B趽��$�׎�\�ko�z���PÆa�����6��j�Q1?(�~kB���Sf�1����·�0�\���82w���E��Z'�9����wGDM���d�0@d*�k�wD�?�ͨU���:�#�<��9R�9Q �<·���a�1�t�"�٦%���Vv�@��#�q�`N`�{l�:���g:�{�� �j��s�۾;u�iMi1��}�w�&�G�ڧ��UƔ��"?ݤ�k�Z\�b��q��O�ۙ����Cy��=~ H�s�xJl#�|�8��j���G�a��ۏ��Y�y�e;�nWA�ؒ������a�H�� �3�����O@_������!N'CC���4�"��>��N們۩�j��=������P�Ĵ&ܿ���@�7A�0�.e�	�ul��N��tH�5�o��]��D�\�����z�F���"R�Rn������̷�(�!+7����B�qP�p�G%��	��DI�����+Š�Qu�r�A?��G��ϕG�����@��=�){W-�s,yT�����F���a,��i����� ��c𩌿�J�<B@;L���;]�B�=6���؈�O�Ŀn͈�{�g�;&
E3��'e〲�(zW��P1 0�Gw�A/0�~�����dʖ9�n{I��3��*|8�����aC^
�W�c�{�W��\���Zv�>u��x�g��=A���J��_�k-g�{<�2S����%������uF��4���wD�"J;
qD���^��ʔ��Ĉ,��+����r��)���# ���	l�\|^b��<l_�p��G���xv��uI0���G���W1}�����~�U=C5%
ԎE�xb�;�{�@����F�N���+P�������Q�p�Z ��Gp�<
"$ ���(p,憑/�\<.���nx���2��xv[�� r�M�O�l���a��V�l/���Q�%�m{3�9
�'	Q�p��g��A�u�J�0�m�7�L���;]}��_e��`�A<	E�0V�5<�m�e,%'��|*eo��wi�N&q����<�)[�j�>4U���%14B� �{K����gճu��Ө�깏ڱ���|��D��=<���q`��$�+�K�G��*�P�
���%'vS�9��T�r����{�=Y{ߋ�:ZX��x�u�l�=O|��iu�� ���#�uBI��h� �)w���?B`g���_{��k�O�?����O�?��/	��$'���r�6�B���'*[��	S1	_H�W�p����������̭�9<�g͗���`��g�I:��I>0ҵ�����m���II�[�dXsss�w�\=#?���մ5�+I$X7�F"~a��C��= �9�^�|г��`"�aq�)��_J��]^^���%�J�
��G�I��,�~���Í��!���U/���Á��k�����-<�R �w�ꪯ�^�Eq;����lB�� x��m�2,��Pn�P����ƽ���gS�
�(VN���G[�f@Ӎc��.����/禃kO5�����׀��jX��k��^��n�[��� �e�r�m��M[Bz���b��f�4�c�Pc�ʶE�n�	0������}D�qsq�+nb�h�$���V�6��0\X1��b氆Q�������B��G*?a��^����#�}����ڂwE8o��6�`V�O5��x4{ ��y��!�<�9�MG47�C�¬A\YXX�z�ڗ�`�Pz�{6�۳��Z�4^��^�-|-�
Fر-�$��	
�O�V|��Ӕ��kxo����!����EC���؋���Ӄ�ۜ]�M��R�b}a���K)�tk��[�����, 4��e��w ���`a���D^�:6	@�2Z)s>��'F�?�﹋}�}�s��}1`/.;�}��m����v�� `r�mїDむ&���m�db=��~4,���pK@t< 7��|�IT�6 _��X�� &��\��@�T��F����t�@ٻ=.LN�� �o�(>ط�շ�fk�
���e��}���?��u$H60��{�nZb	����a`n�Ph;�Mư�
�PD$77�6�!M@.�%�C�+=0v㼿���n �%�|X3��6sVc��hU5��s�H����\۴Ӭ쮾߀�?�n��dC�+u>�t���[�0���n�CĀkz��E�k ��W����Ās0P�m�7�z�FNq��A\Z�Жѫ���p J�lzo+- &�e��l��I���������PnG�I1��Qp��W~;|�o�0�3=,�qf��Ļn����>������L��@>��2������� T�Ye��ݷ��3��эq���2���^;\�.��u��������&��n%m�3L��-b��[?��O�?��7�����DD��'�@a�	#{+��lN�^���s5畇�8Rۨ�H��V������Z�{�̛o�T��(�O�?�����U���R࿧C�Ӱ��M�����ۿ����"(}ٱ��L���m��[~��������Hh�"�Hb������cL�O���|d�U�C�P����Wث����������8��$��ۈ*++spv���ѳ0Y�n���/��	�%P$��]����g�8���f�_ڔ�n�,��uMMM� #�{�ꕐvg�Z���GċU��f�'��O����2��<;��^llт��a�_"��f���H�U���
N�!�*?�:MMM^�7�?��o�����	�''���"VRhTTT]G�U!#� x��]�Ѫp������~:,�5���4zjʢ�
���ax|�j����&��$y��ب��2;֖���(��[����L}�/���O��,��b�#�[����j�;��?�H�� G�־P��t^m�ϩ���i9:ei���KA�/��W�M�T�5��m|���[Ĥa�K�G�_���%�0��#?�Z^�͑N���o[_�4F���= 1%Q��rdH_ڹ�4^-������"�{��6k>�~#(d_t0�=�\q���J�߫���\�{�`�bD}�Z�ϕ���6��W���U��;��3��LS�A�Ah��/����#��Nx?O([q��o�;N#-B�Sj՝g߷o��mja=ϩ����nv�����z�c���4�S��d�.]։	>��od>)Hd�N�>l��v�CY��?3RB��vO������=�'�U*ԃ�/����y��:��p��7�"~pӿ��lȼ�6P�i����eO�j��A�I&���.:���C�m���}��H+��%܊��ܽ�{X��{&��M�O���Ա��_�:z�
%	C�C��7��Nr�}�����jz���)�\[t���,)2�%Z��>���zy����!���L��p��H�}����޿V�����O(+q��]�I{�FM灿�P`V0�p���d�Mɹ�M.=�g��/����?q��K��qu$Ҫ��r��NS�N��ml[��["_8�\x����BDD��������H�'9S��������Q���˙���A�<�T��lE�=<�A��ge)�V�-���!�ba�������>��`���e���Y������
ufef=6׻�!���{�hq-+�)���y�ҳ,��K����^�r*�")^��{�aO���e��{�M����%��̦Zp��L�V��h���~���czY�sa!�@^_E�0���5���X�筝j���ǅEty��V6Jr��߅^��?D����~E�J"��0OX����8���j��s��*׌��K�����Y��}�pG#>:E2Oޜ[J-z�i5���q����)��K�*�����2c�Y�N�:��0�Zv�WSԏ-�b���s-����eK��d�`fB\���7͕5:
z*�yEڹ^;���@��>�0:�ɶ~�g(����u6ɏ�[i��C���	ȯ6jB��1��G]S?I�|�3246�le�yfQ�������s3��g4�6&�r�)��Gl�>/P.Tky3�a���eި�~�]����`>ӄ���/�D�����R��p���.�S"@m��������s��Y'B�r�[ɯ�N��f�L?6Κ������m�8��>m���}��T����h.���WϿɩJ���my��o��X����aS���%]��{����2UЗ����w�uK���{λ2q"K���J�mj�ѓ��2ϖ�����n�feϮ,\���7G���o�%�4k�����1�W+Um�������$r��&�^8�^f�o�@*�:�	����xn�XIr���E:�kQ�[��%���+'�;�bb�_s�"�B�i�;�E�H�uK��
=c\i��x���6>�cr���5�)н���W��Ҡ�&�p�T�f��79l�ĉTI92�+�Y~�{!:5��%�U�q�!�q��Ǜ�ܮ�]?��)���(W]I����A�MV6V�C/�T� �My�9�|nx?�|�B����E�1ݫ�IVC������"(�R����dV~j�+37�jD�t��>=��P�S����E��g�l����!��d2��o@����sT,���=���9����=kde4\ʘ�ض4���*�P�����D�砮��ʪL�T9�q��G��_��d>��ُ�k��X�W��}�ӵ�R4ׯ�}�//}e+0�����\Wq����B=������R����>��&gC���lW7��0!�T�T����E�/b��79^tDrM�|~V:�b�Ϫ�K||q��|�L�n��h49=��n�9�-y�h��u� e�y<�aP��\+�y��l��f�K�I�d��U��w^#�K�g~��TUS���H�%3�����\zʛ������׸�g_�Nv����/W+R���Gĭ8/ie ��u���'o�n>vY�o���b���RN�.����%�4 ����_�t��VV	�[XX/�5�'8Ñ9�w���#�l��r��)���s�c�r��C�3s=��;����
�v��YA?�P��1��*ꋤ��dClxj[�µ;���#���'W�����_:�]�
a�PS���R6�"�9S�ԏ����y+.YI�w$1��[[��w&�j#o�ĸ���S��T)�(o�F�zG�ɉ1$�\�������.UI��Sh�§��
��}Ϊ!X��m���44��B����x�����tiBE��_���/u�X�"ͬ쌀�2_\@5_.,�����W����B�.���Y(���R	[�ū�I.��8�ʅ�H՘��|E��g<Z��:��.ڝWN!��:�(�2S_�R?&��{E��yBε���pzJ�c�{���GuQ�'K3�S��F�^��X�t%z��(O�G��-#1ctǃ��ϝ�.%���[�z��ET����Z^����u��^l啂#T7��ς|�������@�\~��G,��q[�f�M���T��rm�[/XK�_�>--B�w���� ~���^���1�C����������
�;/�v�G��O>1�U�I��i����X���|H�����cl! }���U7�n��9��Q�+��/h�������$���lɮ���c�._��\S�_�%�:?�f �����TuRc��w������s�V!֥�Ҁ��ޑ��6���_?}�y2���Q��BPVdc���v��X��y��s��o��
�'> �>��Y{S�gn�e���.C��-*	�j�K�:��PqV�֦��.��R}Iw���J���4�t�w���!~!����M5����� ͻ�/�$�rm�b�'� �P%����9�4�>�ՠ�c|��۽��QF2��c�w���M�K���w�\�Yb��D�G�l^�ư̙
�":A .��Sٕ�����5��e�~qE�Ȏ��a|}�4���"�6eve_xO�ql��eI������5 ��-���2������-� �s��W8kӺq�0�����m�I�/�s�<�EE�%U��iX�tul��tS��:���ܯ-�5��߼4��Fk�'�����X����dq���0�����1�[)��?:9!=��*W�^T�XP����w��C׊iUA�H�M�X�)rY�G��?q�4��Y
� �s����͍��?x�W��N��Y,T$U��»��/j���Vƹ}.�[<�-�Rja��kmP��6�|��6��O��z*�I�|ζ������þ���C5~ls�~���ϫ����K`��P5LO1I`A�\�\��9����Ǵ�l,��'f ţ��0��=7�^�^]p3�d�O�t�R��P7?�X�z�9f7���dܦ�::���L��P��3Ӽ���Q�qz����6WG�D�.�JR�jc�7�.0�ף��穬�ؒSymG��*i����qd�����ͰX��U
௮T�|��5���t�$	���>?�IhU�˘���p�L�u�
�!��|�?�v����6�oje�v���5��k{�����W8�d�J��X�6ڟ�,�{nx����m}���Jo�"�AQ��R1u�S$JצW #���-[{�Dʁ�#���K�+��Wv����q-~(�V�OtT峥� w�m�z�+ȍ�]:��Ⱦ=��=?���|�q��e��|e�����6���Q��@�Գ��6���� �>�9�w��c�$�Wn�`����Q�X�˳r�:���e�KIs�7�L]i&(����b�x��������FF�$AH���r���[M��)�=��Qy}|��u��8aP7ܑq3r�sh��X�L]nsL�?����]����Y����]z�WƘ:,r��C47�1���	Y�t
~Y.��u��A��8�

� c�dy�Tz� �
{����	ɗQA`MG�4�T9�E=u�G>V�������ZW��G��T�u��"��������/gjV/��(�wWV<�Jd���o��Y�;�u�r���u%�њ+-����P}���Y��z���O|���Q��/W;J͏3u��J,��!���ZF�r��S@����2mQ�c<�����uΫF*h��r�t�Wj�*���m�Q��˧����gV�4O���k��"����{�����Q:�o�NX[f���J�?c�:�*H*��Q*��)K=rr�	��bG(p�{M����i��>P���d^�����:���}EM�-�Mp�z��$��#hګ�+=�G'�i��|�*R�/*�'k~�{#bQa�k�FZM;�^�jr�TИ�z�~M��ˠr��&oq�Y��g�t��EP�/��>Aq!��B��gtq&���y���7%��Bgu�ĸRò����B��T�3���)�I�:[^��=�^w6L@t*��J�Ql$Ֆ��Ω�V]�����y�5�u��^��)��/�+�����fD]2����rFF.�w5�����4�K�|<\����aB~�G���Krc���JrY���7��)�Z���"?�����i����{AG�]й+�U�c\���g,^��{�m�0H�-Y��{�!{V��EWC*����2��a��������	��#�KG�H�,�$����2U�~.
)���K7-2��(^ܔLQ2v�1W�&2T�[�Y�
�]ֹ�ղ�`}���z���ӆG���1E\���Ƽ��𩍡����Q�Ubb{�1�\R���ұ��v6Y�����K7��D:/�,k����]���_J.~w/>�~����=~U�|�8 ���ԭ1g�p>�v$7�o�`G��X���(�/�A�H��[H*�75M�F���~ؼ8x���I�q�5�X�.�р]^��ZDL㶿�#���8p��#@�4����)8����-��c�_V:�������uI������5<��8������ۂ������Q1H��T�#�ʪ�3c�� c�VH9^��X�m�з�R�-���M O\�5s��x�nV$��k/ =Yc���e�&�tB���2�20#�gT҄~����eI �A�6vx�7�䌔���E�hU+��Ѫ��0GDڵ�檻��9#C�#�!��_��ƒ�)Omt�Fpj�P�?9:�-�R���:?Y�y�}�hq�����?��̏�?��_�+�	n�I�J�؟Of���m;�!���c�@3�]�	{(��,{�['���Л��>K�|�G�G��حȭ^�#�X��|q�nd�d�����A�mj]	UX�{CR�mW��>�߱��kQ��j�ͩ���^*M��_X�a���>]��F4<n�B�-HE�)`�'��kH���5��F?z%3����y�Q�����H7�S/kE\�l��"%߮�3�Kï>�d�i)G� jbƃ�y�O �����<���+�(m�7�|o���$%�����Y�5��ṤF=7+�P	�@�.��t�لYOa��%"D!)O*<D3n~� NĦ�D�<`���P^xvX~���;k���sB�CҢU_��J���K*�������.��r?��̓d�:�����ˇ�l!f��:��. ����JK���2g�����FV�O'ЮMP"����ܛ�z�I��[ͅ(�%搨�wԠ�|w[�\�����-�ޔ	��n�>�+��+T=��j�^���?�x�cX�uo���6s��r��/�a��` ��N�@��<���;�0C�Κj�}��}�4�1 ��s�p�|��!�N_<�vs{����/�O��]V8�S.�"�ͧm��Z�rƼ��ſ
��	�6����/�\�Ө�V�s��_k&"��=��z�R�|v�O����\��s���$�c�*f������	�C���΁�R ��|u�(��uۻp=�^�F����/�;ŞQ����Ζ�jC����6M�_=i�1�3�7*f(�t�q
��+�֏\U5��G�����GϜJ�,�'DڟZ/t����PA��kc~�:�_z�jH�5���
��w�V�1�d����ޜ��T�#u��^߬w���|Y<��^�#���
%jR-X���)گ�2��|�'!��^|�]�cz1S���K��Ε�0==�7�C�(�'Y���@N��z7���k��C��R�E!�7!�=f�rR0��d^L�S%K�D�k���t��>*����t�B�����[��WB��k���S�x�1��,�-v<�@D\�J'�0��NPe��YaK��
ٖ74��ӱ�HM��﶑�I ����Z*/R�+��
�+PN��6)QF���_a�R�騖��k�hY3�0��)3~�6�J����t�=ƆL.H�����n��x�61A����N�@4���>�>bHtP�*XmP(4�4���[R���O�6��1�8�W�9�3��l�C#eɜr��ju��ř717�>�Gy��V��C��9�1N ƅ�`fW���Z�-
Lՠ��-� ���H���1��aji"�y0e�
����.��#W�\�4��|���eǐ�%����9q�� �+��Xc�F�IDt�m���V}7qG��q U۫�8��lKα�E��b�i��]e>Ɩ�����M�=Y8���$>Ѵg��X/���W)�?�`Ue��5=�,�)�����{�C����|3�4Nz��ۼh��[���$>n����!�\�ֻ�]��/θ��M ��S}��qw�0��	��Ϡ�?gP_M[ȍ�$�q�5I��̝o&�ˊ�,�.�Z�h_�?F���G*>*����l�(L|��m|c^���I�'Bl5|f������F�E&"n�=l!�h��6����� l��>}������0��U�D�ޔ��l�	���6�m������(���c����Y=�,��~P���:Ġ�4��Y���3���y��ױ1G� 3��nv��gtlvO�I�u��7����ך������%Vl|�����}=��/�u�Ft���ų�M}�+��E$j���80�9�}�����1�߸^�F2�nX�G���UW�C7�̠&�.z(�	�H0<)a�GDMK�u�x�D^�k��^Mv��&Ġb�1�7�j0��Q��?x��/^��x�f>��|R��_FV��u��cb��IMu�2����dc�]E54�t|��쿮,�%�H^�C9����GǄ��3V�V�9#d!�3w�d�`�����cWjW��D!o��y�/��&�M:�vړ�j�ٯ�G9M�l�`ܽX�M����66W.(�#Q6��R�ğ���UF
���QV{޲	�j9Χ�}��V�|V�����

�� s>��נ6U��N辋��Y�����b���O�K�/�*��-��I�	W�����p����!���"t�^�>� �T��?�o+����T$���g��Ⱦ��\-s"O���鉱Hs��SqAT������%�]���8��&����V�d��Kw�`�Ce؍t���o!)ݥ� ���َ�tU�n:�t���z�i���.:_c��#��Lhֵ0������rIм��;�f��D�g!��T�LU
�q���N?6 �H���ڽ��{Ь��~�h��/B�=yV�y),j�����^�Ù���_����^��TG'm���dv�Fs��`��b��D��q����t�%����M�Z��RG�VK�~�S|�\�b7�8����������D3t꒲���R�̐Bۓ�I,��|���Z��o�n�T���
̴xR?���'�Ҙ�40EEB�ょ��;S��8���f\���+9�\�Ko��:gg�<BFz_X_�X�Wx�d�I:�sqq�)���S�����>u�b��l�Y��
Ҽ���lˏ�S�I^�],2�^/��sﻢ�'��"Y�ƕ��>{NN�6�,[|�b��"��/uM@�N/r>*����=�Sq�bW�E�-����O||&0Hc�n�NSC��ϋw̴��2������+L{2�0ޚ�3LZ�����ׇe�Ϥ��S�����	�_��|��J�9����}� ��g]�g�9��nV�f%�"�L�����3r�S�YYY󫕛��#���1j�>3>����L��r�k������^�ۣ�Zʒf�ե��*#|-t#P��o,B�6�S��I�]~�'��аT��5}m�hT;^�Sb��3@�mzP$�OƮW���H�覵�=g���#�zN)�C�X�?����X|�q��ӏw�m$���蚷�q�2Ta�18�pO�F����@}Dz���}R����p�+��!���u�G�"Bo�_�mr��ܷrGf�Nv�d(��s�%-^��JTiT(�t��ڄ���|���P���<�	�Oz���n+FH���{0k1�#"��T�i$��	��p{�z��:�O�*�<P���4��L���p�(���ǉ^�]���_?�Hm,�p�6k	�%�=�Տli�m֋K]��:�$O�d���pr*�� ����
�ɪ}h�K��ƴ���&G'�e��R�n�]��^/L/�s-�"�8��E���op��������Ǜ�P�J{��שʬ[��ǜb��IM�̃�d΋#8Yu/��\6��[�-�������O�xV$Ȥ����-TL��33-�EZ�0�V��R*_s�+��vJ��,��Q�CQ\X������i�G��`�E�}�8B���"����sU��O]V ����ƅ�+�ܲ�my�fk�z��0���҇�N��]�aF)-}}��/s׿3��*%M.]/�זa�B��/F���{-$oW�!���5z�\}R��gC�,�Ơ�G���
�]Kb���8 ����[��{��O��|���o��V�s�aW����P����)�1�^X��¼K"�Z�='I��IǺk��WJ�����9���u��P�񿥌䛑yd�M!�$+#+����#�GFf�����g�P	��pvg;�~�3����ݟu��z�>��s�>�'o}}}����D,�\�r�$��5�d�����7���;˄x���ͼ�u�o̝}�� -"�	�Og��R��rԫE��*�\p��P�e��FI ��g������2[-烵�rUKb���7PS��%.���W����:�qZQ�6?��H5I��D;���-ޏ:P=__�q��`�o�\`I���!�k:9�L�.g���f_g��/����Xt|À��׿62�O�`W�������Lu� �չ�t��K����0kl�����V�:5I�s.KbO�M�3��v�K�'���;���	�MaL��W�jg�E��W?���B��WD�ㅾ�]:z|!r�WgR���@Hs�#�Z���]12]�"��7�	����;�[�]�.��霝E��]q�`:��}���m
[7�����2;S����z��y�K#���n׈6Z����HW�q��xƱ�h[������l�m݌t��5�f&4�2�&�"_�A�O_,n���I�vZ�Y���|y9�+I�'��뉅����(^[mr�x��ժ,�
�z��c��=i�_x�ٵ���`�w��Z����ݐ�W8B�c�{��E��]�(����c���k@�<^�zC1���H�^Q�XF�x�[���rAL�`�^&Q5(�v�zJ���KVw�۵�5~��/����<�-M�z{5Ӱ���3��V���4f�?m8�#DG]��#"CL�q��㙊�3�2�!j^�D�ڥ����o��&�nM�a��1l��g'�{���g����@29��YQ�pt���fY�S)����ɋF�FW����.x�
U���r4�@U���H���W�=��B)/j?�xz��Ç>�:_yQ~AA|�&+	��-[�'�&	�Mb�6��&>���+驚m����K��^G�3��0�A�
��n��̂�.�O�D�{#+�ҹ	���
#?8��4o^d��@�MtT�!κ����>�GA���P	f���E�Z?VI�c�O^�~o�a�T����*:jS�kK��}���#�T��"��M紅%�L�m���9�LJ��%v՝�H*h8�RZ~�,N�x�	�6y�!|�I����{M?uJ=ZmrO�\��g+W�7�T<v�+>�E����Ct�P����`'9fm�5�;%J��2<7��쮤�y�Wvܥ!�kվj�N���̖Y�b��[��p��N��� ֭p��'�tUJL���6U�0K e>��*���WE�W�w��i@W:�"$nŸո�%?Ms�.D�*�H(E1����u:��*+򓯋�N2Tv���X[�]_ߟ;�zC�sB�Ykm�\��snQV�h�v��ոN����d�%=�r3�� ��"�L�g�fzm������j���j��TIש v	���m.߲委$��V֍�>/|I��ybD:^ɷ��p�S����/��Z���@�z��	[ǒ�㩫��7���u�a�θ~�Rf�u �BM���,0I�DΊ˔q�@���\w��w�DO0���GDX�b��x��M5�!�[iqf���W�ʙ�BziI��k�?y-&��~�h�#A�]�19�xmI�H�5��/��,���e�9U�Rq�'L��ׁ�ۻ=��o}�� ,�����)��UOD��D��ߞ8}ٍY�6��֚C\��^:}���K�,s�oH><1���yM~�
;����C���?���Ig'�`�Z?y��7���G��iy�h�غ�|�-�|���p���5���rL����1���޸@o�/�1M:vKx\v���]��hyA�W�/N�Ivѭ����6m�����Bd�ˏ�3�@�z=�M�)�*���L7�w|)�p�������)�td8���ە�\������QK�*f�0��RU[aaB���?� ��>1U.2Y�=��w=�s1O�O�Ǌۄ���Ӡ#��w�/n0�\)?>�}rV��G���xn}���NWkNE�W�K�G+�v���1��qr�m�}�D<8�<��^P��J�v��[?�&�v�'"�~h�UX�o6]�T�1�˪(��FA�p�h��(v�,�?��O�f��߶Nz|�1L���si���s�����TG#Ҟ�����b7�r�H�j���JxU���DzS"�(�+B���}��o,�|_�NS5��[-!SзA�(�K@�-�Ҏ=���+�H���Y�oE�z����SR��Ӱw�{ռ�������]��?����?t]r^Mz(ht�`��~iv-ݾ��b>�(��>�sn�tQ��+�bu�|8�~�q3��7!Tl?�,��7;|��E{� Ц��JC��7 �2���kY ��?�P�s���*(A[�7�J6���7���U�>F��N�p}s���ևz\1���p�+���������~�����}h	�ۢ����*O�<�#G���b>;���0�[椰�ݔR��������S�&Ov��v��M���^�\&��u��5��M<�E��vϝ�U�ԺU��Z~��})�ç��B1��vK)�,�7-P�!�	��aX�;�ѐ�_�&Ϗ��]��ƨ���e�����x��֦~�,�� �X`��T�I���Z�9���͡��Xz٬Wg5���K�`ή_�[���R:�{�J����x�f��fб��pﯼ4�>��ݰ�c=cT[f��v�I}-j��m�w�}���6j`#��n,��w����W��_�C���V/a�Z�*��e�m9��]+�DS):�O�S�7w�_s$G�@��-&��{>i�-+���	�~a��F������*��'}~4_twq�g�>�Mۘfi!e�RSӷ���6e�S�aW��ׯ�F����$Xq1��5�=��ghvpO�h|��Cz�ir�HD���5�V>!B3�����(�D MĹp(I@���sAj���4�c����0=Ф9�n����������D=*�񣐌�p���{��?��j�Cu��ChrpNw�î��P+�4�Эd{/=E}'����]�$�b$$�}��r�!mm��4`Y+�fǁ���T�9�9����0q�#�A�s��|j��o�5�L��DX�g�h�|4O�s	� 6�D� nz���^���l�p����)�*�Tiۼ;[j�V���U�\��,g�d�3��f�h�x���h�/���u���*9�	�~����f��.k�+^&Do�p�[]aÓ���r��]As�K0�݆�1�� �0�ϕbC�= EZ��U�TP���>��+�`X��I�#�����O��(�`EOOB0��R[B4��H���R̢,;� �q[��$�[�*�w�x��p�l�}q@�XW�$3O薊T��Q�:Q���H��7G��i�/i�P���,��$��.�HY\B�ϫ��.��K�����A�hMI��@%�Le�Hcˁ�gH���FaD��5�xJ� u^*bٳie'��dA�cle2Y�Ox
�D�G���w����/�R�<�9�z�=~�9<���D�������4�����®X�n�.��0;�,㶞H���OwR���	/+r[m����S�����tj���l���+�d�ĭ�x��CxG�5�M�p��_2D�H��nxԌ<��K1���v�:��=`����e��d�tʡ�ـT1+J��L^3��3���6��<j�����l,� :�{{�����0��&�P_���s�5OD+ʝg�Zv�K��RMgtP0�� G�}������J�#�!��g��ٽ2\�~4ǽX�09���*}�������T�`��/�@�r:���;��[J��c�Qh,��m��Z���b������ǆ���+����O�k�W��4�m�{S��W}l��������AGMg�����n��e1��r�������.n����h�������FN3Jn�~ �������31��_�xn�n/��0
�D��M��"���iH�J�4��`&���G��|a�ύ�6	�x_��OF����:�Sax��iE�M���sLV&�k/�`QIzW����S��\�3:�'i�8��~�fU���g;(��e>PX����FE(��1��I��ej���y� Y�vG�~�	y�w �FK�����7`�Ps�=�CX��.W"����+�2�%"�,?����nz�.T��']ٝ`"8��I��@�>�?}�R�@���R�hy��ˎ����]��a��S��g3㉵��)�ө�f>�10��X��/��I��/)�d끋�_+*P?��~y�7���{3_N������Jϙ`�2���;0[KK4��g�"�7�o��s�r��� ��?���}68����o�w�=&T���)�?"
n�?�_?�����?P}^�d��P�ԋ���o�����9�{(�SV�#9�f�nt��>����b�M�!1,�rb������1�c��R�0�-��G'v��<��H�/9�DG��T���h�z��&^�y�N������ǭ����	���J�xp^�5gճ��J�R�Q�K�FA"�'���A�ؑ���d|wUﰦ����j�{H���V=�s��n�%-Pݝ�lO���~A�	�����[�[j=�!���ՙL�X{�[C�{ojd�"����|70�sܫ�!b`�̎���n��~���m�QԌ�Dp=�5�:�l��v�Qf/Un��]��W練-�7�c�L� �4y�C �zה�����q�+D���t��<1�?��rs�)�q�ݗa}w?.��4�V��+�����;��f����K���ǝƭy~�l�4�'�K�_}��<�ʫ��=$���du8<	/���/�u�,W�NP[�?v��T�Ӭ�)Ý��fWx
P�]����0�L�5K{�(C�R��'��}}�ɿTa9�PT�5oy�C~~;��u�
"�TuT랍�����.ss���Kt��9����?<�\Rm�8g7��8��zR�ܮ���~���k}���6L�(~֓x���;C�1��Վ�74�3�NsU�F�#���Lvm�ǰ)]]��
����0
���9J�,�r�J�x`f
/�.�ԛ�s���O�`�L���xN*���fe�Z��C����cm�bc�1�M�x�OhQE����ܼϕ!���d�¶��n����Z���(��/;1��RJ��^���MZ3į�Z�,EE38�6���O*��]yZ�UQ���"e>�[G��1���>tcI��?F�el���d���\crn�V��p�|�����7�V#LR_J�מ!�~]���ٰ\��ti���M����"So�F��Hw�	*v����l�|q���j��)���E;��9��?N��t�h���R���)��U�)����Bđt�s�1
7�f��/�����%� C7��O��v؝�e����(�Ԛ�X��>��<�0��&@��\����h�!-]�Z��
vS��)N�>_���:�A$��>7k�3\M)���&񵺵�W[\��tr���f�Wq���W�Mu7�F4�N��"Y>ڬ�%p�������~s;WCea|7��|�t��0��׋��9����m$7����Y��!��S�R�=,#g$�Y��u��a�9��19��b�Z�r�(y���� �t�e��|��3��v��谾8ɬ�6&����n]G�.�N�k�3b
��,~Z�����jR8�yϴ����"�'�Yϳ�/������7��Bl�J��%��C�j���NA���Sʵ��c�����Т�C7g90�w���h�?���˵�8p���7I́?�b���<��Ҿ�J������ F��3�N�3g�0x�����*BspE�J��Mve|B�˦��p�8VFEg�����ѵj��c m~x:�=?����I���lt(Z�k�I�0~�+Wu��}B��OW�J��rQ�JL�|�x�
N�~���A�v��=H���oEE��$S-4"�B7x9#�h�y�*��>_KG�t�p�j�����9�ݚƄ�v;4���N~�E�e��9=���̤*-x<����D�R�o��dޮϾ�?��J�4�SC`f�r6s�	̣¥�S�"�܅�?�Y��#����߫.1��>Rk��F;��O�~uȃ궽�9j4� 1�?�����@��	/��es wۦׂ0�K&J[4ޅ�5�0�ڢ�gEGŗm%J�`?�ed�L~'�U���=�
�CJ��l��)@�s](����ɵP8V˶�L�/��]�]T��
���'Zӟ-�ޞa9�'��Y"	[j���=iOm��ȦQ�����Z�Aw5��y)H��?n�m���~%������m$��/�l�Ը-Q��0A�7��J��l�1	��^vb^ܯ��ce%�/M~�O���/��ZگF�9��bEûu��_�Vٳk��O��(zG�m�׈2{Ș,�5�S_���K�-����w֎�F��YD��54jss�˟A.�n���W�����)�K���������v=/����%��r��7 ������2������Nm�w���Ywn��4����4F�LovY������J�;�	�q!���)̉B���5y��>��C(7��|S��۵CJ��f.�|�4s �6�C�q��o 2���63�VE��no����@����4�a��vT0@䪥�=����2�.2�l]U����֑�	���ޒf��-�|�zk��f��2���Ѩ`IoQ��`=Q!��t�H�u�X�ij�ߥ����7�r��¥�����ƒq<R�	w���'O.��CQ�S��dR�J��� C���6/쓟)��I �|}M��"ƚ����y~4l�bb�d�P�V;�@�`O���P`��d!y�������q�XZ����Rm}n���zQQѿ���	11,taӰ�{'�h{�ׅ6���J��k�+��4eKc�D�]����HT(����aq�W^<�2��X���밊q���+��;uǫ������u�@���N̉4W�M�OG��GF(�L�g�TY�D�-Ou}���d��S�ˤ�ra��[�`ҦQ���V��'�{��)�<nN�G�R}�"�	;=(�182��ü����o��������\E����l�6:�щ\�NqRR"/���4��`\)ڛ�	��r��r��>�)+U��DO}��rJ�>,���Ʋ�������Ly�7�U�ø�⽙���'���{j}����0Zy�V���kUd�.��nV׵��-���ұ�A&}�tZ�o�j]M���㙯2��R��?�]�/~|ow���M^n�&��7yze��"K��o_%�����s_�-��BS4��A�<H�#?,]��7(!�H����
�h��j{�-�Q����Dwˢm}�X[���H^?��	���ݼ���l5ˢ�
�h\=-B2�d�*��B���"@	C��-îXWS"�������w���"��P.��\���Q$R���+��>i�Љɿ!�)<۽����]�r4�KDQ����{=�$�0!�����v�Aֹa��x�[	s1FJ�Vx���烅	0�%�B���/i���� )����R�����N�w����ǡ����Cߊu7)�Ϗ>��i�J�xꊫe���d��J���b$�5>I'���Qb��<(���Z���w%\0����u"8I�f�;��k�ÿNh@�Sw���{|�@PVg16�a�OG�g�(*�(���ϻMD�M�sʝ���9Wm��[��P�?�1�`�ĸ�$�/<򵵠�ր�W��f�<1�����W�y���y�3ԗ���e��=U*�cKVl�,kQlT:ju��H�1��:����J��&�WT"���#���I�]A̓�S����.��;O���Q��9�/��Z��*�VW	�	x��`��S�4V�ɓ�J�l*��p��Q;����ǭ����=AN����׈N�� ѵ
����G�6��>[�*�D�ҵ;�mW�Z�n���!�F.R,:u�d�V��%)�?!�_���ߤ�z��U��R�M�@����n�	�9jqqm��X�}ŶP?�~������e�G>n��sK��x�&�ī���]����)��Sp��
},�����g��Iٷ/qW�G���|�s�Im	v�@��k��|�ōm*�t�%�"�m�����:�������_��ㄿ��'��yUZ��Zoaaո���%zl��:	�1O{hi��'�^�9z9�5V2VDTғ�c��۠�oͤ�+���M�<���=�x0�@M
�t�:��1� �>k�{Z���R�?���Ƴ��P��RU�ȟ�c|��%���#��Β�P~��+^bDE�i�lA?mX:����.u�fE�x�n��qܱm{�m�����#��y�h�ܵ�Y���b	�=�%ޫ�_WpWs�@�~�>n\Q�����R���/�����i����C��[�0ڔJ���Z4Q	B"��[�W�sV�,}=V� �t�9`� bOZ�W���]�D��&�9)aA�,Y��c��\)�2���	֜am_��K�
�ϧ:O|�
r$K��p�c@5����n���4�"�ܜ(�@�cDhQ: �=���ۚ��~̧���G4_�<�8���ۣ�a�'TE� �����,��P�?�"|��>m��6���f�6�usě�"`br�k1V�q���6��f>�wug�D2�n���){��&GU��7�Ş[\�>ͺ�b���jo���/s}q|"K��D4.��������� ΰ���1�� ��o�%p����� �.8��DA�ni\?az��VCdD��Mg��{��e��~��ќ0�y)�JO&q�u�7ϓ�_;�6�E�X5�={�iX�(C�Mw�s�'�[	��8�q�g���Y,�kDSÃ�7P�� u;����Fu���L�6$Pl��Я��5d�1qy�gU��:��{S!���Ӕ�:_����`&�N*�@��ڷ{t���&"Zw2�q$�x^��G�J� �H��튿ݑ �54����!�a��G�.�6�^��Ǚjk��s➹=礻.t��� c�����0���A؝�(����-s�y A������ms�N"�%<�.Y�_������yzpW�0 Jڏ���r�D@��'~l����4�����oMԚZ���[C�B?���D6nD�bޡ�#��݉�R>to������OJ�X)��:
�!���d�b%;���.�+��tX�����|p�`��W����>_��[���w䱾�֒ *���pz�?)�Q)�F�"oD���e|ʘ��OH�q�������FWO�Q��?�W�aj���L�br77\S+a6.97����ܗM��=��X�8���'6��ƺ�Ә��! �DA��4���)�&����:h� �Sk�՜<����}�ω�c��m¨/������ф���F�-�:�{&|�.^�؜���
���{j*��A���TJ��2��zTT�Ep�К��c_E���,��Sň7��0Mߛ�M�+��ܸ�q7��WlҐq_�M��u����r��7rZ߄�׬�lJ��D��N�%�q���?�7��������B�}L	�z��X4ӣ)��tU�,�u�٬�H�̾�<�$<t�k�����Ju'埶�c^;���Բ�M��	��㑃G�	(��l����cƙb>�f��=�i-4:�ە6vj�}�G��Q��{�D��~FQ�(�`�:��9���-�8�G2�QQ�(�}E�Z���W(�\B���M8���τ�	�(HsW�wFl���!���S���0����5+͋+�vU�)�	�~fۍ����3��o����A�`y���.y3���8"B.�u�����Oc���j�mT�Dӯ��^���e��Q�/�d'�����1�*��<���Xa͔��������޸M���[¿&��n��X����x6����l�G�1��q������WC<`f����ܪb~^��S
=���<�W�K�4�B��G��=�r�NQ���O��QSsB��/����m [�צ��h8��Nb�Tq����Ou���o�.����}塎��1$�A$�����GJdaJ�g�;�?s�~�$ɦ�p�=��E�¨i�u��*([��@h��t�3���e�!T�U,�r��e��!@e/�p�W8wY�b:���mf];%%������h��&Q5q�.�[�bE!h<�b}�7;%+�wްE�ޟh����?���ٍ��Z�ފ�� �X-���z��d��S�y�$�>-��(E����a�k�ڑ�\�ٿ��.�ܼ�ܥ:A��~>h%�f�}����%W�ȆK���X�=u~�E�E�5+$�АwRO�z� ��|�!�ux0_��xcҸR�s��S{��Ҟ�3ٱ�)�u'��u(�]���-{apiľ�/K%�e��A���]���xO*����Q�ơ�Ғ��p��N�aV��G@2�ɨ�#�UY�)5`}���]CM��Qy'�Dj$[L.�}uWn�^d�|{��h�����bP�H�q6��~G&e!���D]�Yƽ���7ݒ�ľ�t0�;�ҏ!f��:dW8�*��`�]�s�d�V�#�F�2k��+W���� c\��jh��l��ե�O�&���g�F!x��fga[U�.��:���Ǆ�JvDz������~
�O1���m�]E��P�4#6�t�Ӣes�A�;�����p
:���h4���&ǭW�s��F���YP����!���6�F^�غ�VbĊ�*s%��}��|�0�/Fi��onm���_v:[�f����s5�Kg<+��۪��Mv� ��oZN��wD�h��G�u�����Q���R�VK͉ٓ�m+�{�`�	D��������sT����ծ^����'k��L���[\�����Co�M4 ����^�ZNb�P$�h�ȣ�!i�q�TuZ����0�F�Ą��tq��N/��Ҕ������T��+�|��l��Pޱx
�o�"\+70F�2�n�0	\Ÿ
U~��>Ғ����T)y��JK�Y;,�:|$��K���� �R�Zv�I�Ԍ� ��{w��R/4����7p; ʭͥz�sW�Y��;_H��`�Xs�&���l`�X�	��~��x���a��k�4gn��#�>������{�)�U-��u&]��;P% ���.��_�oFcS�9���g�|t!L�{뀟T7�W�uj^
#Pދ��Е� �Ĭ��$X�s�r&�U���|Z�TQ�86 ��j��E�85Y�	�x�iF:�n�Se���Z��~��Kw��}����ݒ�Ӟ<���OKS����׌?v�������R1nj��?n8�g���T�L�lo�|VthWQ�i�Q��$s����(�ʃYQ��R�>h���	�9�jr�>�F��'uu��~�?r�u�5 f���~B���Q~� PFjn�/#�.@��kA��,�����to���^xV�*w�iSʹ3g�EtM-�j{o��m�]�I��T��*���Z�`��H�-T������`J�)P���s��Z�~��팱�@�?K�m#˻�Ⱥ�̥}-ڦ%�Ϲm�����u��.��������e�V�ꔁ�`�-��:�+w���նЕe
��=UHcG:-���Փ'~{&�A�M�����3�#�n�!��ZS�a��'��k�g(=mqJ��st�*���=�B�I'�y��<}��3{ĥ����5Up�J$_�r]Ȏ���Ums��xR�{ʇ��:U`̡
<�����X��i1��T��1�� %�7���b>8fk��܁�@��:��	�� ����C��t�g1	�2���[Z㮏D�]�p~ry�h�S����n-܂I[\]G�xO&����r�m� ��{L�fi��W���K&���o��I��~��kl������\)���Q�)��̬ۓ���Ug_�6��/!��f�*������@�WV(�^�@���� :]|hpWhF �lr&��kf���pû>ۜ�-�!� 5��̜K��Փ&{���w������/��͕�ܐ�d,YiA���$ :��n۵����Τ �:m��t�M5���A����A�}��s2�{��;��H^�)�O���;~�������E�&X�tX�@��߿��^�(���a�o�[:��L�Jhd'�݄�1T�Mϛ��k�����P��*�F��G����$��y�,+׾�������J���p�Ys���}0����}������ťQ��ҹ���B	�p:�	���>����wiq�5;�`����J������2Q�W�ޯ�ĝ�km�29��B���f5<���]\��J��>8iƯ��]ڷ��3ޣ/۝ ��?�`�'}��G�Ƕ��c�W[�?Z�a$H��V���n��R5���h�G�$l�i�7��kM�-���G�8H��.�/���\n�V���� ��U�ku��6�#Bg+i;^:鲮ii���B&γ;�����r�@���h�N7n��/լ��A�n�-m%i�&o�eB����2�z�ݜ���˚�1�m.�fԬwX���>���cՎ�o�BWBM�@��w�tu�IS�9Z�x�P#�U�۞r�F�v����<|�'��~#�9A\�.х6�կX9� �����V���������m����>�����z� )���FtdQ�{�=9c}������nJDu���ݶ�����d|&�0������)�f�~��!J4#�1G���{_\t�H���]0Ǻd�4AWn`�N�#vl�j��&�Y�+���}���/��|
�*�|��κscT����\�]��x���͹�愙(V �n��Z�Rv���"h��'1�x��ׯ[��zN�l&��"
�٭�͝%��#�i� �X��@�tt����ɾW<�,��>/����\��)�E\���䅳[����U��g����w����b���.E�4�6h�7\����>(���;�����)���9��!ﯠ��`�cS����FY���>������L.ح����[
�bS��/U>��}�|����b�yz�%��w,�����ŝ���;`f��8�e�mz��_EWq�]Y�=._eL�2��S{{�7��	l�6y~�!<��8�}pП��=��x��{�7F9	u����PC�!��f�_>:�5Xx����~����n�/� �%�`���1�	��B��B��N	(X�������2M�^���.��g�q��R�`�y�*Cm�J�7���#�j�f�i|���f�Muk ,��Q+���T-����xN�^YXDF�еFa�Nk'�+�j?ێ������m���������~�]Ή��n_����8	�H����'��^�?��헭��+�n�fb��P�5�������e6����V�v��\����Ǖ@a�Œ�$���t@O�8���[]h���b��Nk�8O쳘��	�=�@��@�8�� ��2(��u����+������8�!� ӫ�$�V$&��*_�&Ҡ�Jfn���N}��� j��m�d�<h��i�B :}}����GJ����ޅ�bm"��Z��$�\*R2ۭi���E Chl0���	qS��x�*��W�n�d:9"))	���A�'�S N���:և�р@�D�����G�K0��[I����w9ܙ�B��*���A��ϼ�-8�W>�z�������~g:�j��H�җ����Z�i�Z�C���C����g���1J�p��t��;�Q0����b2ȟ��Dh��qd���V�?1�����UK���ES�,g�� Xo��8�|{h[�.~s�2&+J��
�ڗl/�£�Wºo`d_0�Ǝ�p^l]��X�����A+�5��K�T���z�ц4VST�nJ�}�m":B.��]m����h!o��R�+�C��>�m��W��8�5j�)�pZW�����=WV2a�+���S��yxxp��85a
wI���k��=o����c�q�&$�NmK�=6:q~`�i���n�_������G$�	2sο�,�j�U���yL�>�	�;�ރH8����=ޏ\Q��������pA��ו!�D�w��{$��n?�ҙ8בD��k���f�o��u##����@��t�N3��e�f��B��� R, G�]���?_�L�ȋ����|\e�:o����ra��
MF���w�� �S�@�Y�4����f����{|��|���-�"

��a�o�C^*V�W�~�ze�^-�-��z+l��'�$�&����g4+8A�����y�0����k@��ބ��Kqq<D��|u��<9GՆ�|�����'"<�/_i�][3�j�-�{�$��s;�N�g����(���]�[������a�������Ҽ޲=v����%/u�7$�pv�
�͈�hr*�8@s�f����Ҏ�@���Z4;cJ��R�}]g�ܔ���Hw����y�f��j~�{����aGW[cÜ��P������'�"{�he�x�M-���A&2���m* ARy[8�	��%Jq��������1J-{a�S��E��<�����z�γmVThq�Ynm�ÊX�V�kĤ��H��3���p���2�fmm=!*��֝Y����j"�����'�3���Xƶj�/��9��Fm�i6�o� 2�*���#�G^ ������K'D�**[���iUZE~�۾bp��� L���B|S�a�v�U�>pL�X5Ӧ��Z2m7�%��b^��y�C_�s:�t���� �L[6G�坝��As�W'�wg��g�@�%��c�5`�B[�T�)��m/����BZ
�=�-<a��ws�,2U��M��mr.�*�0[$�վe;Q�t;��E��B6+��6S}X�����a�å�_FцT;^oF�<D]��X#=^�j�E�"����J��<p>��۠�jH�k���z�h�[����N'K��������A~(*��j�br�RU��~������E@�ҫe%��d�Α�v_ҼL�0�=i��+��
�ִ�R_ I�_��*/75
���C���L#���Ӡ0��_Z�^�l�4.6�9h9��Ӯ+ ��O�yX���0�Wy����LV�,vvv��ee'��_#<m�ȿJ�}��`#��F9y�b��#o^[���J\|[/af��������j�.�sE����m�c��}Q�_�$� �=�~oq�N���1�U�ڷ(j����6��$ޝl-'F��L@�C�U�������?�*g��\v>��k�ɩil���P�:�.�ܾx��W66SYY5e�Et]�!�E���"�}��`�E�3��u����/e���C�0)44;5����N��[2�7�2"n,&�P)K�ƀ���`F���&�D��߲��Fތx���ޭ!�8���'I�����u��&�x5isb�~E�4~�6P���_ѹ*��E�.M����W ��D�ih�	[�^Y�"�]�VK�|ry�Y�}�8���\<0=T6h������f��u-��ef$��u�_n��(4��c9�?�ꆾ��;�≒��~�]�Eb́�n����kC��K~(�w`�j��w�������{�V�@_K�*2��?��8ϒ���|���A另��x�&=�}^iZ� >���ʶ���D���3?4���o K�������̄���~��?� b&���QO	��iB�5�`0�0���*�~5��G��;O����PT&S]�9� p���e�v�"�!:��� 	n�y��p��۫±^?R��,����/��N�n�a:Ƣ�ѳ��� �G1=����Z੖�s%@"T-����Jv�y���Ky(-T��p� ���Q�D�E!��v� �$D*2�2�7g�sUS���G��tKckA��!z������s|3��WoJ}Qs�Y�1��"]��"q��[] ��Unv6��DZ5�i��g��( ���6�|���g#|[��g�G�Z�sl�<�d�VGh+/�ɱh����M��c���%���I�]�N/]��Q:
�^4�e��G����7���dJe�U�E���%6����?�;�qEo���Nh+��Ы`�+��qTb!���ƫ�g���4=�N�&�<�V�h�O���\|Y�VBӅ��E^*����h���PUgdϠ.�ck,�'ΰ������}��n9\��	�l��J��#�0��'��*�8+��k��d�b ^p�Ez��n�2k@d��k�6)�x���ji�5�D��S<-�R�� KK\�� ??R\��/*E�f��ӝi��Ѡ#p r˳35�HV�@�C�n|^�7c!U�Z�y�2+uc�k
����I�H^n�.��5��z���Ƀ�/��NZ����.Ǻ��Db���x�{!f��	d���O���02L��m-�y�mmsiS}w2�|�P�etU���I�W�	�s���=�-��6E%ҰG�5g�����+�yn ����ơ1eWya�/6��_�G C�w�9����v4����v�����	͉�����J�:U�X��F���/���b�_A���8�w��G�=vm�7W�����f.rk�����`���gߚI�w��{a=L�*���E�$�!m����f���ʯ_�*�-|���@R>=���Dh-ͳ�G��"�DxSɶ��e�u���e�8���F��=�ں�'Foo4�ֿH������v���Fp��%���p;�hv��Ή�b1��?g��7T&�j�xe,,�&�����RO ���	 h̧���QM�|���]}���̍�N���;���;���@���q�FܝR��6\�G�Q����^�r|P�ê,m>�g-�@�똇V]]�Ǡ&�*=:N"�k��o�T?��&21?�m:Q>���ץ�+Z�'�C>��MC�!N
@����C&�z}�;���| Xt7������5ա�|�g�b�a݂����O�Gz�L�ÂӁ�3P'6+My�w��"������KH%� ou�k���CH�?Y�Y���S��Po����<�D:�7툅S=p��[�D$�G�e�y����B��4r�x�yD���� �my���ny���;���z�Q�Ɔ�8"�l������eX�N�$l�\�_���~��L�����mc/�;ma�:�s��slYn����p�����^��Uw�,���s�;q�sf90U�����j�+śo���x�US�-����Z3dրzդ=,�,c^�S`��=2��JF$���N#G��cjk^W9����Gg9��s �]I�6�O�S��P�XX�9QR��>�6������:���ޣXV�e�u�_�}u���!��n��O	��
�&�RȼC�d*d+{�D�����v�J${���gƱ��z���=~ޥ�5�����|]��z��goth�.P�U�������W9CK6$i����e��B~���r*<<�4I�U]�ӻ�{�+��Z�0X�K�u�t�?|V�<-���|�d��n����0MC�:wb1��|�و߳�j��|0�ͣ��>'Ϧ�C�����0����?��]��W��"�����N���;��a{U^���e)��Gn/7
Y��a�/n'5&:�θ6돎����g��Yy��A����(�����Z��+m���fĭ� V���ig1�bā��g`4(��;'I�w�l6���	k�T��X��2*e��&���޺W��YM�Zc���_
�#}�,������si/o%IĄ���R��|�Sd����>�3O��V2E9�F}�{<���PǼ���Q�7�g�a&��o�d�Z��ѝm����J����u���	 �롧��Cה`�~�-؜<x�ex�)f0�6n�'���
J�+8��c��E�7���hj��DY$�즨��F��E����;e�t:�\¼Ք��|�r<��S����"C�����i��{��O�v�Oݭ�k���ǕA��=��v�<mY�����ѶQ{K5��~/ӥ
�"÷GG^�x+����i;��.�p�;�����s�>��o�[�n�b��6
r��x&<@O[{�FSf'!��{��0vZ0~
��^�x���?i{���)Kช��+m����y��N8�g Y+w�.s@����}E5T��܃��a6E&�[���״���g��L4���"�ƞ�Xo�EC�Ve�EǷ�$j�n��xH�"=�.�E0�Fk�=�y� +�L���:���z]!Q�j��v�)R�J6�a�
:Փyw]�Z&:q�vE���ݵV �m����l%z��K�[��[�IzX��/��.�����F=]R#l��gW�]�k_]��|+�1Y9j쌇����
���������h�������4�NG9�1�Ԡ;�%�E�b��S%�'0N���7@�M�
;��&�j;��\�;[�X+[H���k�&xC����l������s�CBw~8����C#� ����:�0eϽv4Z�~��!;�Q� �2鞿�h%��Uo�G��kD����k�؎U�4��;
����Mo|���cK��)�I�H��S<����F��W�?ȼxj:4�$,_�|�Ų_`��9� t�Ov(��mH{���ʌ|�.�ҙZ��h�K\�r�(��H��b��� ?;m����2�e�o-��y��3},໊��Љxz���m��=� �5UN%����6}����w
0H�1f�*^��%�@tv'�r&�߱�
`��c�==�I�,�w��9����~I�I�xu���h�׿4�O�R����1��"��U�_��89��^e�ۖ�8�ɕZ��j*8�5/�� ��7��ʰ�	Mh��8�
����\_�]�¤����B����������D �� Yi�pG~�h���Y<JC�/(��)���3��A^�����xD-��[Cxb��-��·�
�c1Z�k	�7/�I��m�K-��%��H�z�o�&.!�73G����(���X��4f����+��!�q6௳�_���%�\U�M_0]h@$�b&{����r�/��B@|������b��&<w�*!��o��
������[�z�wIM��CRpd+������u�6^�$���-�@]d��(�ۓ�������G��A�{v<�`������D�

T7�7�n~�B�`k缽D��ݘ{�6�T)7S������~��5����{�>�'/������/����B��w��ﳓ�8�����RϢ�Kg�$��,.�y|l�
(��W�tA��=E<�+��52e�j���w>g�U����ۋ�\&X�A���� �q�;L.��<V��\̂/�?���@�{�R�x�����Ƣ��bҨVG p�Z[;I��u1�C���7�]/f;��=��H�/�w�@p� ���Hd\9o��e�W}fFY����A͕�g�-���P��_O�����Z�Z��M�IpsX�iX�o�]���� �������y;�Ή�:C��a����{a"����r_k,k���w��_�#�3�Ghʎ��9��Ȭ.�jZ'xNќ,�yh�o7@�|F�?�ӂ�696o0���Vi��s�]�?dTap������ѡ�|y��H�.&�l%�:�W��U�|�aY��o�h0�u��k����S��� ϫ��4��Cщ$�k�ygr�5�x������1~k��:��g��J��d2zs��%�k4'@��Ӯ���Wz;�D#ϟ���p�h�څEz�I�b�� �7��� .<���(�D����;qu�6��K9�*<ڟ/!�λ}�I�v�����������8�DC����D�Te�`�}�u�3�¤�l�@8d�Z���a��z9Y�IV`�u�LN �M���0m$lNrM�������ԇYE��{88�O][9�NZ� ��'_�v $������'C'�2�X���#���BK���������[�Z�[:WS=!M��~q��^���-/80�乁$+�wU@�(�k�7���2U� h�_�̔�~�eG��.�z�A/�)oή����_�I�{}fh�t]�jI�۟p�����Q�]$����P��4�?��4�U�	r���,���uX��Ws�G��Ͱ��'<I��Py����ˣ#��eNa���㮝�����O<	�S[�t������ .*���/����3A$sI�E�'�s#�2���|m3
2q@�;4��y�\mW���T���j �M|sS�I�գ��$0�9�wJZ�����3'�"�3���Щ�=�
4�
	i���/����a��w�ե�f[:\�c�X���Ѷ�3��V�m������m�d��"�X=^]HԽqj���i�)	`��o�)�HLԒ�(�;�<IpU��SwS6"�=�����:n��҉}}>�����~���v?��9Vc)��I�(H���z����8���#�|�c!�lR�i�{�M
x9�� �-3�"���ݭŝ�ʌ�J0����x���7���l,RM�#�H�4�@u��(�
4���᧳��|�h\���OjV�l%��%
�_�N�`���*���o���MjE�h�f��.����c�x@���T�z�'bEOzx��e�d���>�记0z���O����c�P{� ���y[~z���hH�c,2�i��y=**��e�t�����٢O����'5/�m�S�p,l%A��/�P�6#�9 Y�W�.]���ٲ�J���˖����?��Bї��TF�$�q_��W�)xRGr]� �T�jx�*y�׿}s���%�B��ӄN�?QzT=/yQ�ީ�	�l�o4���E�@��)��PV�!,ഠ	�> ����7}`^���f�4=��>�H]�n9�BI�O�ڿ�'Ҳ�<a8�`�B��kb2�]�cQ��qjZ3˼�K�� Y��ev=����)Ӥ��q�����<��-Q&Ў%7�O�_��!oM�"��a/��\�����~���(9.d�YO�`@�`�TM�B��gOv=K�j{C�}�u�e9i{��.9zk�e��՛+^f*���B����ߨ!�����UCG�9�;;N�G�n����^�}w�ttr��&���ww����%�9s>?��J�a��P�7��}4�*67��*BW�*
OEC埝����z?�^Sm�J���;��~_$���M MQ@�?�N%W���fJ��qA�� gVZ��0����7<I��t\W>�c�(ē���t�*�5�������߃�a�LK����W]������������h��q�q�ؠ�ʜ����`z�Y��{���W!0c��.�#<]N���h =�	�6��|���z���V`���G��%B�H.}Ar��.�J���r!��c�A�62��ʮ*�L.Vr��q6SD+�1�Β!2�C��\�� j��}�Wm�I����w6�(��c.��t�w��S�9�4�=�s=#�IvK_������r4���뿎LZ��B�[��e�U��5>��}��*O��&�Y*U
^\����g�~����SHQvvBU����X��ګ���N��R�J���m�D|�9h�ڀE^��W���0�V�����'@��Z?��f�ǒ�/Ah�'�$���lo��@���N/TM��?��$<��fjʚpWr�w��嘗 2 ��g������?��ub?�#٘\����ܲ#�_�B�bOD0:Dx��~�Ю��2�@�8K�;��kyzzU�e�W��"���2���{}�L��^�2N�
�k��� �&�<��x���TD�=�*�q�S^�2\~����\��|+�8'#��Ht˿������Ơ�h��A3�԰�P]ِp����Ç_罥r��R�u�q�s�Ȫ��DO�~ih���%��!��և���A�ܜ� ������앆�"���g�#�T-���5�^�<����~�+r���I�|}X���Ճ�/�D�<�<���\}�����Ͼ5ۋ\eG;���jhkg�H}=�l"Mv�b�
]��c�k���I������}��QC5�A3���+��h�=�?����fRn��ۖj�WuUEE˥S	��M����Lѹ3�>'��E�<����}��e��[B62Sk��!m�ݳ%Zj�Ꜩ�܇��W�~���a���6Ž��oX�-�(�Q�mh^�!������6/<���a�q�0S��φ�K
�a�-��εn�!�7�-���4���s�/\�d{��u���o��-���|�X�O�h�����c�O�(��q�v���D���
$h�sE�+̦�Yh�ưY��v0�������~�?˩P�u����5�Ј�
J�Ru;b̥�j|y6
���QG)��;?l�(E0]FG�RW����e�x��2v^`&z.[B�������<�0��#�c҂��n��2�/��]����A�CFJt�p��:1�	U胝�"��n�`�r	30U?e�9�F��$�smw��ۋ�9ą���{��Ч�GAM�+sc�érr�����d���	�{	de����h�;�ĖG	��"�=�h�=	��X�Nݲy}�?O�ͅ%�G��I�t�����ش�9�G�W��XGD���qC�l��8�~<�i��D�<�dt���x� @��g[c�o èȐ�����K��C��ǈ���;B�8V�,�/�-�]��b�|Ę����ߘ��S�sO����0����}��q�Mf�5L8̩�ǃz�L��]f L�~i�o�����M0}�楝�DAk)������N��q`\�+������`j~�p��V��a��vǔ���6�!)Q�Q�(��m'%����S�>_�vV�m(D���^2�h����{��菑���ю�b��:%힟ҥ�����M³�����L��L�Қ4IU�`3�����u�E0�x���F�Ĵ����!����~E�6}|��[�l)B"
NYY�����`F+�����`�iM���E։Q�����)Mx|�<�y3Aۉ���i;��I�"Z��8�\_@�mj�M�r�y��/L�+R�B���,
+�����ׅ�?��+"���]�:T"���uhY��\�E��K��'~}��R���g�?�列M����鱱S�$>���d4����V�}�ť4�o0�M\D��5j�x	�ӏ;ʙ}��XR��7��|����|q\�Z����+�Dz�x�#}*��ئ~��s�m���~��\�?/x�@Ѿ���bH�ozx�f��a{���I���1�7"s���� 9��'�ͣ�	������/�C��1�`2�_j6���Tʦ��s��g�/�����$!S�h��ϲ��ܑ��I�3�-PF����w�p�����lm~7SD�
�#> �*�F-�Y

�b�廖I6L��՘���Yo�M5��qU���
�9̪ �\�dz�Lv�8���VR��B=yigH��V��H�Jb�ױ�hMLT�RiA��=�WNR��]�Y	��o1��R4�_�?h^��nrˏ5y3����
PSS�,T�-㉋6����piޗI�H��YQ�U������L�S��g��D�F��~\�2..����s���l��\Ǹ��ZB(�Q��#��H�H<3ǉǡi��f�(N���ڽ�B����Oo�5���百�q���'�C���?ӡ��3�v�CEL{��!y�+E�n0c�F���}�܈7}g���^A4��=BK�%�[��p�&P����@��������y�ȕ#1P�ϞE�j�p�lBy4�l���k�U���4>�M{�E��ٻ�@�����<�cǢ��enm���?2���p���!翱\U,�7��D�3!}�t@늸���I���mrO��'
��φ|y��ҁ�ᛐ�Ԥu�D��V�7�����|L�+m��?����ׯ�a&E-{�����7��7SL�Ow��M?���U7�}�j���CY�����sJD�;�@o���S���e����G��z��6�fq><b4��������=��:����fv������9��S�	�����桡�2Yf�i�P<��W���\ɳۻ?K?c�f�b�x��̢'pB�az����O��1����p����Y��a۲LF��#�}�����3��=�2;!=���曈Ϳ��vSqr ��oӐ��,Z�����r�S�@�6<|��pne����R��ؽ�>���g&�||��T\�F���rȻ���f�u��f�q��oT���Qm�O|c:7��C��c��1&u�;>�B�_��XVPME"	�W�|Lg��;ۣ��䬩�]�����ѧJ)�Dz���Yu������������ve���{	�K�*�y̤s�?���{�m[>}~�^.���)��7�O�$�	��?@�D���>�k���]8�+ Q뼆��O�0S�th=�������U/��,�fgZq��p%��Bo�S��,_��cõ��|b������˃?��)%f�J7����V�n�<c�Ŝ0�cCÎ���t'�Q�v��cm�mI/0�D]N�x�ң�OyS��ei�!�Tf��;�e���;k���Q H4%�~u��Ls���p�=�wL���8i�;�N�;J�k]�=[� �ed��Pq���d ã������Qvv��I隢U��#K��BL�Tn�ƽ��]�,���ز�"/��ol��S`������pIo����L P����/�D�|- !Q(r�X��B<���'J�pjw��rq�ه���"��<��;aV��?�2�:����
)�I XN���}��M�֛ŒxY��//ʪ=v����<�1�u!�*泺�s%��M��]G�7��������:y�
p���f�P�j]8b\H��#�-��T�ъe��Љ"kF���v���ϟ?Q!��� y�^��[�iJ�tK�"3)���n	)���(\unH��9�:]��i�m��8fY�#�,R��3�����<�R����<n�F��������vq}w�5��[�:��~b�{�$4M���XT�4���L��ad��Z&J�+���������Q7ɴ�UB;�`��I���6-�� ���Д���'έw1냊���L���;��FY��k��3e�41��"�r��'�M�X����!����w�2��Ը�v�
O��������@rT�����̜�ޕ����mg-�����������#������+�m����>cb-�H&�$mц@s��*'
B'J���s��E����LL���Nt�:Lɯ3O�cn�',���RY���V2v6�.��_bn�"A4�7�rTi�A��c99t����Y�H|�*j�Z[���x𷫧�8�]Y�*��UfF�ke�����Ky��ػ^�к#�1!�=�1�>ӛ$�N�|����{^{�&"�E���L�6us�;��˭kř�6#��>t�N�H��׀�V̑�u����Zq���{S��ȇ���f3��X^�U�r����.h~aAJ$Y�{��;c���]M�abe�4rH��_MF� ���hD0®?��\'=�H)<��f[���F^_�Vg�ϙ�Z��3����MnA��������I��lU�L&ߩ����͓z5*H�g{;��4�g����Au->��/#��5��M���OWX>����w��iD��MS����vI���-бۭN�����!5����B(�Om��Ji���G�j+ɽ_�m&����_���W��gqr��w�2?��9B2�>���H[ɧ|��Fѡ�x�C�vp'�i��pY?I��<c��;�k���K��VV8�Ct�C�?�3��w۶��B��<�o�	����T�b�`RFu�46T�,�V�y%)�Δ�ׁ�H��H�����4�dEσ�`�����!�R�ݨ��R�>K���}�0������\�Ȉl��>!�w�*��0q&�rzz���,�
pN&���g�R��&�Q�I�L"��k�@������'�����	YF|��~3/ �/�(vZ|D���@{Y��ф�m��z���;&ʪ����+1E���5�؁@�����ٝa���VV�t�|m���e��p���LunM�h�f�N���ozy�*)5���Ϡ�;Z{�ի|�6��jH�A-�V�G�88q�(ܷ���)9a��]>��왅7G t,�g%(l�f���u`����r�M]��|ORqs{�HS��k4 u�V�{}��q� j�1�5�G{�#����h�A��7@�?B��Xf�3�ƈ��,+� ����ǯur��0a76�|��4���s��oO'F�$J3ݮ[�P����Үk����ߚ�,u��̶T��d����Clu�-Jr�"M~9�z��>E�k̿x�tt���H`w���O�9pc:Ɋ|��A�ڋu�����q����h�����C=�bՎ2�~I��i�|fѼ0��9a#r�h1g)�b�,IUu�.�;9�.��� &,{Y�]�n� �dnn�4�"�1�}9j�� ]H~����/��uM�{K�u��v�[$�SS?����#Ζ���ݣ��"������`�2��
��^7�E�Ǳ�2&��+"�%ɯ�� N��w����l�LC7li���E� �<�Ln,.�z1�ޅ�A���:8΋uWtX��������g6>��<`bGg�|���i�?��}��mZ�L�0?i�X)ȍ!������a����}D+�ߍ.��}<gX1!�޼�Y�S�	ҡ?w�������L}����O�3���
�՜N�&ڌC뚪/�3�[�B�����Lv�X�9�싛%ŊNak7�3��dO��\�v�+Z� �w��>������4Q�d�=SNa��7�"˅� �4]��ץ��dU���� �aG�����n�V�⣂�J�Jk(@$,��z��q544t����1�
%�A\��H~�&�?���1��x�����EFizϾ`-r�+e=�Ą+�uO�rtc�*]qM�G�;�L������Q�GF��޸�P�SY���S��v�0���1���o��d0|+� ��ʯ@� ��އ!V6;�[��������_��,zFPR�x����E�i>�����Ҋ�@�Lŗ"��[=�}dTuJ)x/�Z7� �����!��9,��)ה��X����/ 6�dLxq�֣�f |�bb�{��h��W�khp���#u���}���$��y��1�ID�mL�3���" a��B��.����󾋵�P���DR��VR�.*`Q��:��@���)���q;��y��o�Ÿ�#�+����z����P��1�~R��K���KyEK���� 7�����M������X�D6;�ܘ^��}��_�[7��y�-Q1�	F������>�Q���+W�ca��2��{��h�����(J�w���k:�*�DA��zuZ+���&ex�$!���w�LL�n/���7����_���2��� ���b/e��Mbẘ�d�$Y��y3�$a�<:1;H��z�xҌ��~49;� �x�Vk�"��D+x��cG͗��	�@�%]�d��XK;vݛ�Ρ e}K�А�\7��X ��$��?[~&��d8T#tg��K�B-'��4�w)��LE��SN�L��ő�*�T +���Q���(F��&��k�\�}�β��Z���ּ�d쿶��<�ϝ/x���TC��1�y�j��Eu��=��i(KK���DdB�[0�o��??贾4,��X�ޅ�(�L�69��-`��+au�+͉I�I%"�ƂB��(A.���5u���r��j�ƗT�짼_���;�2ln��)�(�����Xk=f�@�*jʘ�H�c�T�N8�pD��4��	���6�=�E��\�\ ��D�<C��<�NA`5\
|�\T�73�	`3yv�HCү��y�){-�.Ud���N���/��\rF�\z�y�3�0i���k��"=iD�C���g�W������CD{�./�A�q��Cu�	O�� ���?ѿ�TҤ8l���jO�����\���� �s$��/6��V�E��#��5�;w�@�RU��`�$)�������� U�bn˧'�c��s�p�B�!�U�F8�j|��B�*X���}��L��YF-��!���<4��ነ�T��^��X�j�R�nq��*� B���Ǟ��U/�e����^ �8:�o�u��y6���?�*�gm����A��j.�����a�j�[[?���8�4��gѻ|��s_���i|����a��/c����~�|��1~#��ǘ�A�+�� 
2�Aq��M�ӭ%� ��l"Tx!������	d�Rs�Gm��@.khhhY-�!4?J�[�^�n���̍�7fݚ�����*��E��ѹ1��w5�˾^::�����ë���R@,-���Ξ(��OA>6�ީL�z*)�~7o<G;�b��)�C����L�	ɉ�^V �n�t��Ƌ�_�� �Z��繥�	:�:�4�&Aap�TR�F+A�sZ��pSu}+�w-ALU�`�qz��`����'�V�<����=����.�g�ݺ ?Q��/k��`e��V��A B�\�|�ҝN(�G m�it*��&4����<u�������mW�)���E����]��Mov�c͞/�C5f�
(~�ƶ�w9���w�!�1�N��$lR�lx�#.s}Ӛ�H�$��\c�������*��2�����VL�L|;�`���G�@J�JX����bw�d�w,� ��n��}KO�r6z�V<^�q��@�&���1x�3BK��!��YF{��3��Z
��Z�2����a�E��O�m��QA�N����#Ǚ�*T�;���	�IL�b�`w�� +���e5�!��[���G�|,>z#�zq5p�W�<ZM__�SRQ�C::9Y4妜F�� �Q����z�ve$������-L+=q�|y�5r����_�M���j�~��A#��),_�^0 9�����N��oې��L�s����B�U��H�q��dYRu�7̎M������<�ݯ�
\�V�U �Lw�E�T�JN�i'��Eۇ�������ba�1W*�B�>{�&f�ѹ�������}@Y{k���@�ܺ�p���D�W�/e�w�J��B��@�����I�][{e�~-���)|�bC��e�3�9q�F<Hs�nm���<�t׹��a)��ѫ�:t�e�{�_^K*Qʒ�����h����=�ݗ��e�������>=�t�fdtRS�[�E�틮ʁ@��J�|�5�=-��OX��L��)t��u��u�{��ؗYO�x�Z���j�����3K�e-�gjo�I�SĤ�=-�z ��?��3!�dwNl`���=��Q���ȳ
��s/��W.)�-,�E,�q�Y�z6�H1��*jw�V{�jx,�W��d,Lww|�n���O�����k���y>��PYm[8矬����'O�X߷~aq�^z�6�z��/�M�r���0�����%���7�(�7�4}S�iI��Hn���x�S�P�A�An�*��!�$|�<x;I貌���a�5�{K��H���^XO��H�O=�kv/Íb�,���#�}0�t�2�J���� C������;�(���4Ϋ�v�LUS%��"��T�&H��s�o:��R>��Fa\��TqRqA���Jr��_==��,\���N� r�����
B�ɗ��G̒�C���Y��U�U����0H�E�6�0��R��ʽ�Y��^�fq�])s�5v!�����"h�;:��waBdXh�laՎ��g�I��'%Q�E �<^�'�󛹁�f֋O��y�%/� �M�߬�e�_���2kc�����s��̅��y�:�_�%�6��Տ�NqZ�4��&�j�yE����%��<pL����lx3�5F$ �����N:J�%�zw=���텿�ο/P|�Y8�U?�jkk���	3�O������l���D�l�R��&����qD˽�'[DJ�j�9�$���U�-����;`�8Iq1�#���3����a�q� d�����j��^������_�L�����a5@������$⧍�b�?{���!�[���#�l�Q+mQᥥ����9̒�x���G�U�8�}9SB<����_9���� �%`�� ���{��ͯ ��Cnإ�W�V>��bm�w�����NChғ���qm���) ��ٷ7����-��`c��P_2��k�b_�Ր��k*��O�s����s�ʸU�'k��Qv|� ��D���I+��I�U�c���w�����]�j��`���Qm��7�4����(Ғ��'�6�8�T&��s&�{�M��z��ԧ���Nr�99�Ǻe ;�}������.A�H���ibݴ��7�-Q�&� $[w
5�L������� I�ჼ�}Ӱ��a���%V��[����_�`pc����d@���=����W�_VY�U��V�&�Ĭ�Q>|�q�.�QwÃH�ˍ�':01M w��ٻ�t�F��ِ�$��yL��<�	�N㪩���I՛�R[�1�22WvG�ڜ�K�]#�T�;�<�������e���i;s��۪�{KÄ��mH:m�"�H��k��z����wݹD�`�ὅ�
��V,�z�F����.v���d�L.��/p�[ZJ?x���Td��&+�(!����ȯϊ����z<���mҝ"�R�jm�oK7���ou�L�hp���r�������%C�?���S����oB�R��p��ަ;*m{�U����o���.U:n��v�Lr�1��dk����c�+W(�+���?�b��dd��-bbb[S���XT^�%`�L!�6�6U����A~/���=�⢽Փ��n�9�'H` �{:�S,�b8͈������z]s�s�%��y��f��f�X.��r�T�V�8$�>�%#�IB����>�yY��hU��;�S[�q�����/��R^I/#ϭ0��c�i�k�[����Ƭ�*��p����s��N_�Z�x��R��s��Ј�nq,�1�M'�e�g����}�pzү6�4@8!I�(����ؘw�oڧ����C���HO��I���s���EK��W�����ǆ��ߥǓ�d������HPB7o7A�}�VL���|��CLL򡬠-��x���y�P�0"�NqR Q:̛���6��d5��z���f���Ҫ𼆼�#���Z��� �-y���#��ӳ�7z�tSX�n�r���[G>�H��������7+�hO_��^��F��s!8�c)
�y������Ĵa�~rHG(�iJl��;!�'�F+��ӯ@��7��#��\)���OkB����:�H��9��B%$���l��.\�LE$�c��D��sJ7�+kEh���;8�-\��id�m/�]��L��0�ޱ����ߘ��`͉�)��w��R���B���e�.�!W}��v�~3�*gS�M-�+<��U�S҇�p����]��`g�SFO�^��ln��Y�3�㣃��k���>J+��X���A;����>�e�)�M�#�����QʜY�y�n����ا�0������;bl'�m�d���v�Z.w���έ�7u�|+'��?�:��Aw��6V��:�*������S��VK2/�c�N,ָ�R�ߗ��(��O�|u؞��"߀�s������A������:�����\Z�ZK0��X��w�?�������z#Q�6� � ���.�z u:�޳��ddjbbtͭ�Yo�&��2�&�f�k��Z�l̻{g�@D
r���b=�(3���:�u汚ged�@׎ȇ�t�I�AL3�1 ���l)\�е��y�yY�!���	�������sJ	�c��]�ѣ���TP ���{NIW����)��2LIyy�lw�٭w*���b_���~)�����?͗����3e�v$�-��%,�}�j���	�nB���C#�x��
VZ�f�YEu����tth ��d4�U����!�ۅ��W �D2Q�\���sn�T]n!;K]׫7�+QS+�6�
�C����[.r�O�!�?���u�Zj�4��\�1�`S����Bӯ�������-��8��O<�@���s�I�k��H�s�	iu;]8��D#���C�A�E�1i�I�-m�Y�M��G!Y?x�E�	�o5������}�7�BC����|f���I���9{EFf�?�|�+/��H+,Ru�R��d��F��)�FD���B��7/ ��Z���ri��>;��#�߈4���������G\�x��țs��7O�W����5�O��*7S����/�BV��]B����˻BB�ᗆW�ɘ�e�<9i���u:������7�k�����L�-�Xq��Y�t�[ϒ��}	������+B^���Ks���v�Ae@u�$a��Y����_g<�m;v1�T}h빮<B<�:�;��Xd�����0�� H�h���@ >�=Uut䥤���tr���+{����;�p� 11b�g�)$Y�XP:��ajSm�6�ϋg����yc�.�D���m�l^3���`!p}2�����̪�>��4z��=}�����H��Q��?�#'��u�S�)�mL~x��n�J�����w��6A�H#^��$�L��O�Ve�S�1��v|X��EjPp��[�[r��'O�(	��*����S����gI
��xGr�`i���^�����|�^�����b�W�j̫�	�֛`^Ku��D��\�f���"�!h6�5Q�<k�5�VV �>bY�I������.P)]^��x'�Ġ�#�ڰ�(u^W��K�/�A���B��/�M���N���b�Uw�OG%�+.~SLՉ����X����ƢB8fg�W㡀x��ׯS�E[.�WF+�}���傸��]`��4ȷm�վ�I7����,��<�ƐY�Q0�gcZ?���8�?�_�N�� ����)�#YeAη���ppp8=��/2�m��r�hoc�y-M2�e�n�^��۷���01�M2Q8�E�fs�؁��}���ip��xks��mx6�pz!hSP�[\k�b�xFo�V����Q�ɿ`�A;9�B
dy���� ��~M��{�o߾-�6R$h;������K\�Q�(�ڃ�M~(Cu
����3��4�YW�ߝ��wsމ�?Xm��M73��
hI�)1Ƃ��Σ�����P�՜�Ȗ'��3���;c�����j����}�Q]#��[�4���0ژ�E �:���������A�'t���FAp��]����j'�n����Se媭�G'�fyR�/!.vHiP��C�Р�J$�CB�jʧ��ɑ����Xǫ�ƋIܺ���Z �7KK����*W72���M2��澗�v��Vt��������:=���qތb�srhY��b����h�����������i��}/G��׏�
�Q��O�
������4�E���]�day���P1?�I�xO�x�u��0j?��ޒ��tz!�Ƶ��l����mS�Q�~�P�:����7$@8D|��i� ���_64�*0ȭE_o�8��%n����������Ɲ�%�Zg���x˻Ȣ�1C�����k+��v���Y��DDd$�����ك`,,z:/�j���2KzPS������.vv�V.���|� ��]�?��_�'�U(7��:#�T�����P�4�
333k��}��ק�A'Wȵ��b�E�����te���X�']A��3��Q�껶PU+�Q/T `�
����1wtvJ��@��[YA��L޿)�O�/��죝�b�����At�;�,cL~U�,�NK��9�U�S��nh��T}�2�|[O�?�oC3�
����t�I�CZi0ii�ƃ�V/�r\��5ر:r�����������U�M)B����ث�%���&3�^=���^59���xbw�2oeeX@�[�[�G��F���V�1孒�wT�<R�����}�_�5=��W�{[=��@��~!Y�b�}�j��I̧��Aش�QZ�{m�m��NT�"Eײtɑ������b�/?��o` �N�B0i��y%e��%��R��V��, �Z��
�ӛ����M
E��?a�%j+;�L`J*��.\.����Ve�
���`��?������&��$å��;��S�h��D�;
����?��g����KM&�8AsRp���En#Yߚfg��%1��D�+e�"�m��
�������0�������̷���&�ȡ���(��R
�)�O+�t�r��y���u�9%	'= �\��W L5�P� ��G}V쎱����	tNT-dp���͍Y0�6��ջ��4]�1]�W�M�hM�����%��LP6-���"O��07w��+s�?�^�n;�WUo �4iU��9���o�{���e��	��`�IE�/��W��,����^�U�`����򌌵u��*1,u������rK!_����s�T���,��h[%5�.�Vh�Ԁ��9�V �����xJN0Ձ����qqZ���a9�i�ٹ����)O!�uJ�C1f���z8���f�#�z��[GuVt<[<^y4�|+E��'��0O	�^�m�`�pR\�	�J7�����F_j�r�Gl�<j;֣������d��)�p&I��̦ũV���uݳ�%�A��$)�������b!��RS�"���~X�1��j�Ile�� �zTde����6/�Hc�Olt��{��x0u�#�NR����58Go?nF��:˭��}-Y�
�bŷ`-_�6 7�����N�MA eUTh�aA�������wK�W(LUɼ�Ng�?i�I�p>6[���J{g��� <�;�XFmk3w�j�/Mc\\�}H7�춼�,�~�:/���̏�ˣ�v��s �kbЉxKa�x��P�s�B#���ҧ�(~�tϻSz����)|K��i���{(`q"a=ڔ�)G�44��S�Rf';���
�>��#N	Xߜ�paN<��Q๏�C��A���z
)�X!/y�	䪇3[�՜BOw�_���!Ȝ��\xe"XV76p{���_-�%uKݡ��Z���� GLc���q��ơ۝��4�q���B���P����pQO�����K@���� ��;�!�={�����+���jV�#I�t� j�Z�8Q�-�R�@��R3��BQxC����j��lܑtxb�̠r72�q�V�1<�&��rJ�=��ԓFL��v�q0�w���Z�Wo�־�������Q�%�Q��VQ@���PDPR���.���DBrF����]���{�_��׾�u_q�5�AO�91O�7�r��3�MT���� �
3�o���_�!7<�u�1�ڗ�B�?��_�_�k P���s��e�[c
x!�-A���d�����k���
�ei@VFu�G������߿Y���7�V��	��O�+��nlQ�����@?��c��]�!�o�ٕ�V��˅&{%��#Ne8hLp�7</�p�'t��\���z��F�޼;����,}9'p���W������^�[�R̹g@��;S����[�
L�)~��hڗAf���9�_z�WLz�ڈNN~>ٝ;w ⯕5�
*C� �~��`�����낙��+�H��l����!6������͵YR�@����v�/��@#FRR���LU ���	;�f�����5�d��ds*M�GY���Y��9�[4��g�,��Q�0�
�(���wApj���ͧ'ީQЩ���Zz{��d���@{HKKϏ��{���@�sZ��&�k+s��v�<��1L#<�\VWH����A->D5�g���m�I6�]@k����׭�'�c�J+U���Ѿ(���a��n@˵�<߮�6OM��u�>�-W_��C�����v1�٦i1ز7�V8�s��oC����d�]�u��� o�g3��79O��l*Tf���#�g;��۹�s
�3�	
�}�**�� Ki��@r�}p�;D�Æ1�R�5o��{���]'H��1`ßJ��#3(�:�I������K�rq��;�(33����7ɥ����]	��o����ϳ$��
��)�o �������?(�_5�,�,74�q����'��P�A�7׷�yG��.�8(�fM���b||��kW6��y�v���y�ovF;�1��!l^?0{�.��	�Q^��>�]�z��O[1F���pkjj>t����h�d9���bH�L��ok����.���O�nO�c����Q߹V�6
���� ���69��w�/MT���FV�>|��t����Nݽy����Q�D���d���Я�T\���i�C8���W��vm;�b�Z������H'4��E�Ӎg'�i#�m��k,������p� 1-�; �<@Y�,	��}F���R撛�٬9������C/1�͸CG�-�7W��omi�_���f�#1.F��,�������{���[K�7s[{��w4Y�e��{4Ѷ�>��:�m���菱�)��5.\N�'}9~�ή�p�s�nA�6����w����h�q/�L�����k�eCnOz�PE��n~z3����8P�=B��c_�]/�3���6qv�>��ɭ[y��8�n�/����3(�`�!*������zR\a�A���A��9�>r+��$��������Lb�&��Z��B�X�Uk�ʯ혱s��zGV[˦`��%�h�!�._�d�M�|�BW.tU#p�!S�_L�R��ʪ��k����(����n	e}�/�����m3�5�C
�9�bRF�|�S:Q&�`6d����GS2��T�8��Ӎ��BG�|�V�0�il�����Ϡ'��\ �CJH��� �[�������;��$�ۂ�I��te�GW䦤/�ɜ��p�?}�,��^ֹ��������(��HW�8���3���'�������g����5 ��OS�ƽ�x`EBGG�KC#<����E|J�i)�k�������Zw{��#��+�m}�7�)��=.g�a5�ܟ[s�Z���������g���1����[9?�ᶂ��ۙF\��q����1����Tq���A���W��lD���d{�����8��Z^>�W�n>�##_55�^�Q�F�Mi��e&��#�m1@�g!�M|=w�2�&_��Ńg�'߯��Q4�`w��8���私�I��������v�|a�v��y��;n���d4���rO`������ĩ3�y� ��հ��u׷�:[�
u���I��t�@�i�h�||n� �_�(�p��T�g�@��(��o^�
J
��/�?c��WU�ի9����9��Ƈ�� �>Ϩ~�����؂cbO�R�Y�4x���=~'�x�*yk;��u]����>���w$c�q� �M�ܰS0���e��I�#�(]"�6Td���ݠ���#=e��2�m�z�2<o��{��wZ<�d�?y㌛[ZU���+]ԿcL����w.w����v<X����]2:/5#��ۣ���9�L(�Q$�Kz��,R^F��n��p��� ����ULu��`��:!1��c/��P�A�Р�@�/�ɑc� >#��t�G@D�e���SL�MX�g��ā��À��Q��I����<��D����"�Zf'�z�_��~0�S����$���|ږ��B�W�$�t�Xu�b�j�]�6�,���.�Hs8�#��J�����w4w_�I ���s�KC�/��w��Ԑ\��N��,SE��z�,�e��8���U3d�J�gj�-I^�jgR�w�
�wr*�M�c�"޿#�[t�G�C���j�}����Nh���H����z�ݼM����֜��?�Ġ�&oC P[�6�.� �����5V��444B�*Ny{^�7�pz�M({�����3���n��RD�隭x5[>r���9�Dz0���1��2�j��c�4m���ǯۗ?�{�x��֩bU�=���I�x�񳫕{��}��,�Pe��9��PH�B��5��;����A}��o��}o\���y�?����R�]�ckX�����{j��4�gV����."�ա{^z�P���Ⱦ�Jn-�k�_����5K��<����ٛL��_|��9}���dLgZT�����c'��rt�#�#ȁ�_B-����&��4&��O��w���M�$����Q��}�ժe7�z\1z�[52�tMG<����4?�5/���N��=��ٓ�l��j�E�3Rl�Ԣ/�#�Ɔ�Y�5��v�����B�@�`�R�*�bS��m�c;����=
���QY�6��i�P����b�[��6[3��+ȁ�zO�a�a��U����KGq=�Z����ֶm��j�Yk �=�S�����.�7XhK��u��"|l��X2:��x*ŸxAs+��ˤ%�������w��u��Y�`V��R��l0��6�	�x��s�$�G�Q;��3�v���6��kc+���o�:�������[QNfY/�S`�:+�>*�c�>���D'�n�����cP/��"h���#/�����(��DE|�_�R&ɲL;3�.*Sg�ί#�]���g��8�94E��d�_� �|@��(Gg��!K�ծO����b��-��G��߂��Lþu�2n�0��z� '�k}�*/D#�B?ն�_&�ޣ�vb&�h�BoI,Ѩ���u�%�/Z��=2�c�
���]�����Hq�[��pV�F2�"tSC�w��}�f��*�e=�2ϼ���~���N|fR}*���mjG��rK����)�UAx���/��*t�Z%���M�{�u�-�'�*��˼��7/�]u��犬Tee��uP	��F�tMJ���X����ǧ�m#S-��X����f��!�7��n�<�Q�4N.;X�>(�Ӗ�%�Q��zc0����S��/�0����n�[Ld�����N-���c�z���0��Ɋ#����!�5������vo����~�����R�*�,�m��]ak�s�+D2>0Ƀ��|���,bv0EŊ�)��̫a)�B��җ����HV�����~�Pϴ �bdt�.m˥C���;��8���_�#ð�9B���d�!�M��/��]�h��._9B�}�k�p�A�lAEy	��#%K2�Ը�J��+b�j��� �r8x`�Y��zOw'I�wq˙-H8��ׯPQ��{�wv���f��t0�9�3�O��b�O�
a����J5�fj�F����QMmY��W�/��늻$bD���Aa��M�4���I�	�����E��.�FI�#s�c}0%�̀9�o
;ԋ��Z��P�����}�N�۠�#��	�E�т�)�#�[o{�zކܝ��5�sUl�=���;���ᗉz+����IW�%BtW�M퀔?���SU��9Q1��а�-�x��J `�je;Z����)�t%�ړ���h�*�mc����ϸ*"Ilw��H�ڹTr�'
����9�敘�9-��9ڔ���Ixf�~�T�V:�_��b7��:0�V�l5ߢ�3��N�7i:b0wM�x��zC�����K��%��v�B���OgPq�E]	B�@-��N�h����8��U�{���ܠp��ޙ��R!t���-���M1��Nһ-D���]�ajPv��=�һV��1� �qM�����r�#Vā6lr>6??��@�9��oJ��g���Bޕ
1L5S�æ���z���=]�۰M��uH��1�������Gc�
��_�8aLG�O�T�$g>� =����-q�b�a�C�_1F�$5�&�t
���E -����*t��/�H�]�d�&ǔK��SP��Y]��A�4݅B�����v��
��'JC�Ĥح3�zK�Du_���ճ.��	�P��=����:�)�Om��������I�����d��y+oX��&2�}�B�l���)Ѥ�o�K�N{;��Q����}?�����<#wZA�i�ua���U�F��ٸe~�yw�_rB����/6���2��C���qE��o�ү�]�J��/B�!��j�L��\\��g^Ӿ����g�/M1�.ӌ�̰�Ł��G̼뗺 �n��
�:^�`0�G�R\V	��ș��L}�љ����hvq����/ھ���"�
̤�4�ba �p&6ż�K�Q���G�3b���
O����r�/�W"܂�,�0��h!bH��Mb�C�B4i���e�պ�,�a�_��^|bK|�$�*��ɾ��"4�	��^ 4+��(<�M�F�1{Ok�z��}��.$f�$�A�/b��/�=�F�XI@�#_�����������˹��-�f��*��BG�N,�����b��:����X��>��c)0m9���<�����^Y����S�����9	�ТP�^&%m���|zxi{TEv�WڗXW�(�|ɱᎿ���c$t�N���h��+����i#S�n_�h��m��[g6P"	o$��!^�w<�RH���Z��X�G+�^���8�d �<�\N;�8c�hMo�&��/�p���4_��
j;$u��@y5B���(hs�����J*���P�(f�*�)�)x~�hu��ڇ6B R@0A7��&r`�Te�"(�ET��Z�oU�t�Dy�COu���Y��~Z��y��a��%F���s�H���y}m�3ֵ���wT���{�&N��}ϔ���mj*�r�K~�qH��\ѧ���z� �g�{��N ~�rz�ֈ@��S?]]]1u�z���8�L �n��ZrP�nԶ�.�'�:oY���А��1$&~/ �չI�w���J;���]+8�=��;�.��wF��~L��~�8J�|�9&����~@�d�$�' ��Z���Xm�D��V҉9}�}�QpH�M�C72F#D5���c'2�X?]���`*�YgDp�K���$G	��f��"�t�!c�cu���.0�d����&_5k�x]��X����]��헙�x@��u5ಂ��A	�CD*��;�Y�8�sY��:�N�Ns���'�����0�;R�Q)��l�'ʫ��)�#�ܥ`��Զ>��з���e������2��g�h#6�SN�e�:���I@�S�赧�5km�QS��������>PK6R[����?��T��9d�����a��-�uQε`��ӡK<R��qN ������c���)~^Ow��3�W����췂<v�s@�d+���f���"�8h�8�I�dY�f8@ɢ�!+��, ��� \)��yj)���twh^�q�!,.%z�zΔ�h7��4�L0�,cɶC
�ҳN���a�� L��~���\���tl$I8��w��/�1J��_�B��PoN�݅�Wx9��B�0�b�Y��z�r�@=��\��9�c
fTtc<�=�;��,����9y%��n�*.�+�ĩ#�:k�U��`wB��є�� Y�To&KGi�G�=��2�R����;�+L�"ppX�%p�΋O�; NJ߬>�p�����ۿ�HxO�k1K�zn������5K�"�.�M�$>m�HNF�C7RQ�mGoqa���e�D�7Л�?{�N��di�m�_�3����੻
��~�ȡ���L�斛z!'�N��Qu��v��{q��D/�����`�+��_�/Wc�U'wA��j��9Ze������*/XU#��2�)�a�i�!`#T��ż��ВQ5��O,��~>@��Y��@1�E��������pw�']/��pU�=��t,ƾ�X����y�n���7�)�M$r��1����LP�riIs������{QQQ���.����bMq����MU'��+3ܖ�zT��qy�	�[�wN�;����<�zj����b�a҂��2Z���1��$�?dpH�yeg@ʩ3�f�����Ϟea��H�IN+.�JM����[;h��� $�Ē�8�Y������� ���LG���/��X����^�I�YFl����W힞a$�y���Z��9���zo;���%Ơ�?�h;��L��N2�k����lw���( QH�7�Z�+�x �^��E4[�q'��2�,����أ���Y�����.����b����1"������f��U"�W'Z+6����ʩ��eX���R>�h���'���i�i�f�f/7w��d�1��"J� ���XOKQG*�E�^��i5�o% v<�1+l����{��.siQ;C�GR]O$�訧��	>�=,0;;��zY ��<�3޶@>cm��e�r��7�,Jl����<V�G�s��3ܕ�f��p|�B���%�ȯ�>�����>1N���^�U�B󭱷[�P)�f��5����[ӫ�l=9Y�x^ՏDې���$2��A�B ������眳y�LK۳�0�/vG�rw�4:""�pcmT� ������q�&���=�A��s��9�m�����O0�VgŸ��Е���L�*���jFa�A�P��lyc��pM�y���N�h����Fr���\���y*���U�=I��/7\��|�%���م"�G����/Wuu���;s��Cz�ĀfbC�@��"�b $�X_�a�d� ��;�E�p�"ߗn���"����L�W5S���y�{ܡ�3h����?�j{��eu�
n��\��
�:1�T�o<�C%� )�.\�外��w���c��ʬ�G4��<w��Y|�"	\6 �R���bi��+e�9�9�<�y�V� $d1�4om�m�"�gq��t�K��SvJ�����n�?ύ��1=	wl~	r
�1C�ٖ���-��"2���\�n�!"hpre��i�:)����͵8���T!w�^�#h��U�V��F�肦mыB#l?�n���4;����a0�dQz{�Ɇ�y�-�M��`�;��\�R�_��[����2�`K@ctN@����uD���A*2\�rI��w@�>{�����s
C�Xn)���'��7zR�Wax��"���9��Q�k#��T#�%�0�h<��K��tpV��)��*�@D�O�g�6F�s��f�}~Yz��l*Q�+L>��k��ELO�[e��d{ =�Y���&YN��x�*�%��9��7�!�/.�k"L�itc��������ߌm��X�2퓾?�U!�Cj#o��i����� ��>G3�N.�0]��n[��~��9��}0��O#qq��+���4^��OW�R[{���'�g�s� nf�ƈP��A�X ��rl}���:=�/�=L}
T�T��,3>�#u��j�=�a�i`�)%zD)F���-����P��!�l+t��F��FzN���Dn�%��R��M�I���X������~���v�6C�&܂���5+��+F�8�N��n�O
~����z ��^(
vl��~,!^����6��ޮ�=���)H=¾b$.89�7*�ԙor��B��ީ��0}7C�M&?۲�*���Y��8:]��c�*-5) R6�)�n�Ϋ�f�)�,ae��O>����DV뭯'�#���:E�C��Ŭ�]�������]i�湾�8�Yǽ��Wr�� ��gq�C`���d54s���	r.�G��͇%���N�����-�|3n��p�1�J[����- Q��E��z@(J�-��%�m:Zփ�f�K�M��E�nف(��yI�N����8�
I][��>SWWw�{uB'H��"A����(L���4��s��~��'�Fd�٠�$�����k���O�1#vKU�?��A��Q)y� �Jފhߝ���Ӌ���iN-D2�?ߴB������u����@�+�|S�rWw��r�*��'l�+඼'����X`�l�X��Zo[�*3=��ɴI@��0��1��ah������*V<g�7�E'�N=�[���'^�f(M���C���|,��Y�l�Ȏ�W���h-�,���"�[^?o�f����M|�Ix5�b*X>�dժ�*���dKH��q��ΝS���_�Hq� ܥ��҈�mм��75�;�&|�d�sk��#�y� �өs�y�YM4�����=��@^
�䥢��&0�U��lI=e�È�|�?�	D�/�h���B1zj��E~E���i�Jj���Fu�2�=B�0A��l�������y$e�H
��Ƴ�2���U�*mCL���!�w=�c������ʸ	��������pQ�����S����˱y�D�5>��g�H�M��,��1旖���x�W��*�hR/�<p%f�-����ì����s;���Ҝ��aQ�R�,�M��˛r��YdJݡՆ��{��;��Ѽ&~���[c��J��灼'f�A'�����֭�4TXC-&ߛh��4�gQ��P�0�&w��*�1eI�@�#��9���n%!1j��/|&͕.�r���`����<�7))�ܳ<+tj��Ol��L�iC7KI%bD�W��1�a�M�@ki�1��ͽ��#-��ٜLqsz_oۤR�ʯ��)�J���D��#�^�fEp3ۛ�WU������9�y���p������<i�6��GH�c^�+��I��[\��>OI�7�R[�i:V��3���s� ��m^s+a*���jJk|�u:5���]󰠱E����}�_�wFl����m��Xa���xσݎJ@＇Բ|	�"�9ؿ�����ۀ�dh4/��G,�ϸ����"�G�����n�4�ٯ�Y��H	��z���W�?�8Z-�`
l�������~�υ�t��-c�6�a`O7FU������K���x)����t�M��)'}��nO~[G�)�!�n�qC��Fk���wT����'?�ϲ��t� ����?��o����w��Z���[�S%7�_��t��i�Ͷ{Ov.�ϴZ6:��vJ*�M��sDT���T�K�//�;L���c�G�dM��g�-YcA�\[i0.�ِ Uά�v�����Z�׽#�XZZ�ZG�$T�^O���!o�O��=��N��M�I�"ڶ�!YVH�������ta�T�Eܝ��&÷��N切������.��/t�F�\��η�*JKg	�n(�̎��G���#��������w������*q_���wY�&y����s�z⛽Qۣ���7̬��s��9\9Z$���<���C������
A��q��O�{��Ӎ�y�~nԮ�N�>���!"�~nu��x�s�d�UQ�ѯ�
\R����g��6�%l��l����p��55�\�H�O�R���=���I_DĦ)���?���s�Gc��*�`���v8��|�7�uA�i%�G*{eأe��Y�>־=�L�EAM�N�9W��5$x�ط���D�"+&u �3>�Mz�N�~���Ӽ��,�����Rm�<M�T,;��8�O0Yf��ꝫ�~�/c�(M�k�=�i�r����+t?SsS[@y��0�n��?�i` ���A#C�{�����E���Z�_o:�;�\Q�_�	)��(�x[x���R~��(ByH�`�j��ZE'E�S,�;��x�~(�V����e��1���@
['kmx���L}�P��;���A��а�a#�i�c����bgF1����1��5�Gl�L��&�t�u:�R&���m�g��G� ػ�*��B���)*���8���4�ǽ(?�`���T_�*0 ��7�����0�����g1�XY��ʇ��+j(�����d��D���Y�A��W�ґ�z�Zo�n�{Q���cJ*b����0�#�Z>D��m᜛���tT��re�\z �.�u�q3�Qөy{�9V~��iNh�Kw���X��R?�tä�z�F掷��~�pɝ��}�u���c�J:�1�壟�T6�Sx�8����-҃��T§�`W�8G���n ŒԆ��5�E/��iֿ��;�C��d����{l�tT�ak�"U��U���wT�޹]�`�:�wiN�����2%7���rU$���c ���Yni�ǕL6�?����(H
 ��f��䦆�5?���I�%���9:V�2g'��nv�4�i�L�t�Z���3C�}��=ť�6�2�[m��0r˫�+�.�>�p��RX�V�*;��eZb��>���n�����K���L�.9±B
�)Óe��W`xZ[�`�E=�F��}T���*We����	�I]�}$���ɶR&���� u3D�&l�r�L�R�"�6�U�E	U��Pqb}��q��!����(�Dew����8|m-�A�tM6����w��U���<��䩏��f٫\�̕ܥ����aѵ��C�Q$�ߺՔ�c��Cl���GMwe���u���Ċ��}��O^���7�J[�K@�X#��1��|h�ba��}��uh[�,F@k�m�8U���� ��S�~P*h����ҹJG�؉$��8JD#�X����n{�� ")4��\�'����y{`�ͨFfbw��s����i��3K�VǛ���_�����tS;�����5ox�8����՗���
��Э�3�;ƾ�RO"4q)|��<u3��L�2���A �ˢ��/��S�NǲE�j�/HO��$�E=Ф� ��W��K�4�W��leM�v��S���?����:2��_�~��>�.��}��)$��h��Y]�X�Z[�@ؾ��
��M��6�8~��s�ERF�,�v�X7�;b�`�������}���漪Un�������o�`D�6����im������>5e� ܝv�Ï��b�BЌ����7��$]ԣf��֨�d�i%�_�G�k��#o$2͕`d��Zoꈪ�`���Hz>xQ&p=����R���n64����l��BQ���f�`�(��^�h^k<i�(J�onH����ĊX?_k�����;��H ��1g�_��{ah�U����% ��R����;ȶ_A^-�t-|��N�;tq,o��.�h�Ѹr����C|���_�&~�Yr^�)N��_�{#����N��5�ķ���2@>��2C�7R�T'�|S��L�EI�x�g��"8 vn׳��ҕ�f���H�����δҝ�9���g��!��\|d��ӗ^�Zș����tu�:�d�#l�4x˹,�7_����~ ֻ�h�TG�%�"������pYɴL�X�Z�~�H��z�Jt���d�o��6����}�6���F�* ǇZ�X?���-a�w�^F����k#���G�L'!B�Cӵ��h=B��v^[�'�B��M�4]��|��T*�f
n��}c*�/7�v������%�@9L�~(�*b�&���3q0u���!�.�ma�񽤤$����g��	��G=��g��F󐒥�I�	g�>f���DK��@Ӡo[�4��-�;6?g�uf[&_/�n�� W�0��t X_��ڳ4u�_0���8����*ܸ+vaaǉ9]82��)c����.���A/�	�ǁ�m��wT3���if2{�};
���{��Rp<�{��6G6rUf^i��BT����7| ��/T������^G����H��[LZ\����)�j$�G�1��WH�m-�"���1ZP>��dՇE�RL�|�������}��b�EMR
���}�*a�ݦ���:Q��sϮ���4�ͯ��lfG<�K;�Z�#sl�O�y��fv��"�l���tŧ�O/;-�������Dk(K��M��g-����`�a��{'w�(��}�6�][`-rt⮚�� @���4f�a��Y�ۖ�%�]>��C��^�4S5��y�Ax�YaL���?�*v���Au��q��XrTII��N�y ,��yF5������A�[���C�&��/}|�����L�Q��a��DTxU��k*��ц���u'u��P'3��t)V'��q5N8�K-P$&N������$QS16�h�Sy>���_J���A��'ن�b��p���$ˏ�k�p@_tŋ"�s@w��;�h�+����$A%N��"	�s�(����)��fx���O����$���C�bI�i[�Wv<�4�����6,�#nu�K�&o{�a��o\��ba�=^"�P��#k�G=���&���"�?`E��*����D�w_���]y�a����S)��&\����4uy��Y��3"�V��C���y�#L6Hv�-�` ��W�.%�(����A�r��[�i�]7'&Z�u*i7�g�����CN�hZ�s��uC%z��w�W�W�^ea}|�6ʑ�7��g
�,�Z�mj��5BR%Ε�h�W�N{R�d��P0d��p;'-�I*D�\)�.�
�#��I�Wf"μ�QUr���*nxp��Cz��	�@Z�~��)������J�v��
5g��d��3Dbne=���1 ����Y���1bX#=)��,����j;�'�T�@��NhGe<
�q�3v�T�6l'Ȝ�x�����n�����Ys M���/`������A�?HƣN%X!9��ԧ�C�,�&�0�8�͕�ۢ���㲚�S�`�A�x��:�j::ox-R�kMS�|
1Fȩ�=�5��4r��+&/^n�@���YM�a^�.h"c�5"!�@S_X�q�f2fskk^V�6=BH~�؜������j��hRm������|5st�4�P`�j\�;�of9�V�\l@��������<�*i�Y����w�T�3���K�ٸk�[�m���v��p�I*9��<���Î���_�7�D� W�Ml�ܶ��ߠ������l��ۊ^��Mw�dT:̈fڥ�>�9sr��v\��X]�N�!9˯����Y1���y~�Ѥ�1Yi�M�cR���L*ʥv��C� >)�
1g.��e��v���^��|�|��*�D�tW�O����:�����%���Q����5Ҳ��;�&3e���	�������,�Tj�Yw���HL�r˦�ĉ6�^�L�����Ͱ.��F'v;:�;ׁ����x���ϩ��k�?BR>�54�z�T�X��V�/��]o�d�\�|W�ǨLνC�i%�k#y���4@�4�<��z����j��[wŊ����Y�V?�ǅ�|b���G8�.���лq9L����M��g��"o��ŧ�'�O{�N��%�ؤ��v"�#鈦H܅ΰ�m�;=�V*�>�|���7쁹��ۜ��q%�}����� �9iU�F@��U*Д�p�y��f���C��ԇU]0iƨ�!���؇q�1"Z�t3��c�6��ku�l��	4	�3Ύ�S'�wu�E�l\�_�\|2���M-�����ϛ'w`n�A���t�v?S�#e(õ�.#\(�2O�RWlV��ZO' �LB$���ӧ��px�  <�f(��C���s7\	�QPЦ�u�c`5c��N�?h��g,���I��Q� L��d~˸/
�v�8�3��X	'ggQ6��<�,��c��ςRc�'-`�i�{����=[�k`�H^��k� T`$>�,�dUI���+2�6��%747QJ��6�%��W�7���9����~g8�:�Μ� -㲻49���A@��
攼�
��������J�������j!	H�ɷ��G�q?�ĈȐ2���@m��U9~h��^��S~���hg�<'�����? '���ui����%�f�ܬ���5���T�;3��̈%�����P�:x���ɝ��˴�ļO��P����-K#cc2��)j�� :G��6�������K�{U �CF[�D�ǭ��<G����rVBL�"!�}�������,-�z̖KϠ+�ۣ0I	��Gj������\eV����J����Ƕ%d���R�7W���Sx�i�{��� /����6�_	9�KF�+���*��S�A+O[1.J�.9��p@��q���=�14��"�,�w��6���U7Kn�N�r����x#_���A)����ol��,/ ����$h��O����-��At�	Ǯ���1k��x�hj�wĲ��n�V����BS��$J�n�r�l��?t���S���<�9Z�,Q��)��ިv��6=�@.�eraS����t��[���;,���P��f��<�E���D�D�S�?��"�\��/�<9%ڠ�2������_�<�-��`���� ��U��6i^�V�𛵕�N'2y~rn�s���te~%�O��Ǯ�fӕ���Nur_*� ,�š��C)�l��.n�6^D�aZ�6�"Va�t�)%)Tjꚓ���F�*2D�v�U�9���6|�
���<������(LAE��S�� ��◫������rC��;҃QS� ��G�l�����>�!������]{a��9<4҆�tT������y�A�a�Z�on�ˡ�_��[�`0�_��Q@bh{�� �Ҧ`ǟŸ}��>6��+и�zS��i��x+h��ߒ��m!;�,^ECƮs%�R4������?�%��)y��X�_3ӛ�F/����������qPa���X{��KST~�y�6�dR�I_u��WDRY|]"#~�R֮>�:Q;g?�#�k��w̷��R�CY��!�y��ڥB�#�f��7��̻|=�G�������?��%e��z���J���Py�:���1�C���E�]e��A3�c|��䪆\�r6�S!eIB�j)�@���[JR����|�?e�]�!��U�y[��x��xma�	"�+�r,�+*��n�����i�A�ct#B��d�b��ԃ�ʪfcW`�K�7^v���;�.6�=ʧX��\ �F�ť[��Օ{��l�3��؛��sk�>��:��/E�1`��f��2�Xː��@W.���0}B�vژ�F�� ?�^�4����g���u�'�#�"��J^N�ħwh���A��b�%|�7k^�$U��f������
�O(���|�m�(�8�4�_��k�̂�����ee�ޑ�&`#�I��� �fl*)0�Y5�j���	��.�a�WD`�������$��=7��Z�=_�=����]���%?e�;v�w��dP��gA�Ci�>���'���A��[�][:���Zj���s�=�oy��m���{���P/$�$�t��ǻ��2�QW�����䗛K6�BB���<��8���8�`��^u�]�g1gߴXC���&�r��E�����w���%��3�` �=��0x��X��!H]��v����K$0x�i"ϰ�@����T�+�x7'J{��6����{b����? ybٵ��sH���c�����ry����w���М0�g�)U�ˎ3f�@G��{g�ew�y"k�����O��'%M�\��ck�@�'���v�I��_�!w�xȖў����W���s��5a������Ì���~�O�o�$}ek{ۉe:wòZ[�ʯ��.����ٹ2Ϳ�*��#����y/3:u1t�f��x܃�'�	8Qz�K��~>7�Z���\�M_�/E_�X�$���(r���³Ĝ��]NNNq�G[o��L����
�`rJwܝ
�X{���,�
!Ԗ\���^c|�a���I�wA�����nN ��U��׋#"�֙ØDE�+07�F�����1�Y�)*�u�C�dK���OYl�0�.�䲏8� e�����p�����n�`	\&"�S�un��9�d��yc�p��s�'F[�¾W�Ҝ��1�����k�;���S1�AK[ '��M#��dS�f�?�Z�|{vv�VlZ����W�v�ʼ��ua��7�P!�f�)O_bj����'�D�'j������?����#�Em1u눻x�ݶf���|#��Z#�r���|/��܏�S��G��.:K�+I������Z4��'`U��"�U�a�?�b<� ?���	�U(B�H~�˖sE�dk|�]d�� �� u�kF��ٍ?��+����*=nH�YVO?�I/̸��!z���?���.��Oƾ=��mWF?�{ȸ!�<O>0��O�8��ޥ�H�:�7@���2����5���G�]|��rg'��@�8�"lM��Pi�@z��j��(G���<�H&S������( �@:"-�33��,��I����ew4�4�<sa�uk=j�<�7;*Ѹ<�z�& �ތt��O�C��m2ŉ �6]���S�L:��$�zt��&��?m�ş��ֵ|�}jll<�"ml+��9��|ᆴ|?�+�c�8�_k�ȅ�ZB�WF?�<���5 �,O{��PCǠQꨶ,nD�2z����5l�-��̼1��)rt�X5$L�V~����qU�}��g.H�?�"A��ㅗ[ܤ���Lơ (���W��z�/��t��-od��#���ϩ���2���7�İa�uw�q��h���F���^lh�u�ݚ<�a��&ұ�*���Ւy�8'�#��ԣ���y��D���l�>�PWӬ`ȑtY��9vH+�W��Ǐ	�n.mӉ��,����A�^� ��]�Q"!1�/�t^���r"C��
�Tr�}jSa�c5\��(��֣��/��U�����z�qx�Mf�au����vvOQ�T��E�Ĳ��HBb���p����������y�c���s]�5��7�W�Y����t�Q�o���e�PfY����ԯ�E��ƶX,���y[UDL��mp����)jW�\GT�D�C��0i��[K�NG%�=dNI
`O�0!qk2D ���AS�r*�Ģ�c�w!��r�,}��!���n]�����)��g1J�҄�j\~7Z�g �[��yPd
y��f���7Ta����D� ��J*�Y��-�{}�+T�M�Q��w�@��fdp�1=�t��8y-��@��%Y� ���^�y�
�##%u�o]�IҾڊz ����z"�a"B��\ܺE�R!���=]�@KUU��R�[��Tm��(X@T@)*UPi�U�������NE�� E�  ���;����(%@���	��y�w���W8ə�ٳ�Zk��9dqY�̇z�tI?�;�]?w�1z}��%�O��-��['��o
^[+5#�d�Lf5I��	�J�*�_�����`�'8����l�0�f�#�߽�|8f�}y�+��82�bU��8HZ���E���	��Z� 4�4�A�Tb�7Z��3��<WA��gW3}�V�ng�[�v=7<����7�j�7������Yw��S�&�t�	���h�t�<+�>�%(��[U��#�s��y��Z���$�Z�ANV��rr�,�
b�9g��+��;��=ɘ?�v�Ur�����U8G�n�R��*�,��>Y�&#`TYX������Gk���c��s+�X�=���F'��S��hg/�Wޣ�tז��*l��ۭ�N���UWVT���*u�2��!���-x���t�=���� g������c�[o�\sQJq:TS������]2K�f���+�;,G뼢]�j����|��`�[
����������"UwHe����r`�i�����nU&F�k'k
����Z�Z+l�
�l�}E��������� �W�����@s��r/�̫fL�74a[ �"�*e�(B��R4Ӎ�6 �Yd��)3P1ݙ��^����SP7H������qAk��p�Ú4����~Y��_��S���[O���Cտnx��e	cB�$�o=�\ܑ$�r����	�� rы���R1�"����Oz�W�O�����7pw O���O�J�]5:�.����AF�ȴO�b��2o3��8Ŷ(��o~�+?�?��t�y�P;o�={�k��Ub�6K���}u��)0�뱣v8��ڴy�B�a��;/X�瀔u���R���q�4�6�D�;�'��t��B+������SJN�ǣ�1��u�� d���Q3qZ>�R/�{����iIܸ�Y����=�m�R�$��j�^T�ħ��坽݄l���Ë�7N|��|�Ea[,ձO�6�y�Qo���� ��7�~�<A���	��O5�_ҝ�Xy��Ç�k60d5r��<��|�dU�n�r�C/~�C�u���w��m�HC{u����9�4���R~�u�����g�VH���a�N]�~6����8�����s�m��#L�<9֩	&C��',�����v���V�/	u��Gu�#�a�6�[���k��O����ʡ2�Q��3bU?��G�W
)�U%E�w�L�6c�5us�g�ь���9c>\���uk�"'#�{q���5��ʴ�rJ}0��Hu@��Q%h��Lˆ���I:���'�)%��o\&F���x�y�;d������'W(�ˆ�{1�`�
CJ�<u�EX��$ڣ�)c�CYAZ�cAq ���P&�=��Tm��4�ȟ� ,�D�(zӂ�٘�u���R0r:��bG�f��5��@cZZ�n��/��КEWJ���>S8	ڎG���c�w5��	V:����ZOJ�L��I��C�����]�x'=Vg՝�}�;�c��kK������q[��KXz_y��F�f��4D\nri���)O��ʆ`�̆>B#��M?�FA�v�E��lh;�v�;��\TQU�%0��\b�8()�cп�<�5��Ϟ�z�bX�N��{��3�;V��l��D+��Z�b�7
E�Ծ�N&��7 �\�l���X�(��X1��FF��6��(�����_�~�2}��O۱�rOΩ���"�}�u:T����LV���5�w�'�;$�����$��?�W���Ÿ����F�h���f�6��M��ՏgY��'�r�(�S�s	�r�P��P$�S�Sm�l>-zwy* �%V��"R�	�������>[CM�vK�w|3��h�&��8��|G����k�Ć[ę�j�r���.h�Zf�y	����0�>=��H���Ky�Q�q�**�<}vK��H@�.�v�j���2�/�*ȝ�RW��O
�me�Z�&�"�<���)�J"?�)8��ů�o��f�Ɉ<g��6��Wi+1�I��	�싏m&�*y���b;92|�s��T� g���5Z&��a��g,a��a�\fkP]�����W闼�Iͻ��@�����!u1ɻ�~�o���Q+5Pa�����rA����#K'�y�o/H�n28��U��J�h��V�.	=HL #�_jq2�O���	��b�È��fw�O,�v<��-T��:�]�e{/�_���f�ݥ��7��퍾�?K �i:\�gv�C�ꇻ�hըv1z�͞{A�=;؈o��������K�g_মT�5Ǻv|�+���ԘI�R������K�0���c&���P�-��?pB	!� 9���Ȣ���ç4�\v��8�A��"_ʿ��H��b���^�I���w�^�}��8��443�arR��66�6`�����#��\����NkG	�0�Z<�)�y�S�M��� �_�2z6\�s� ��R�=�C����6�j?l�k<��r�%�Q����e��.��O�қ7lp��G�c�Z�m^�kT���v;4N͛��j�j�����Ⱦ �LLLH#�8>� 9i����FxG�zj�E��V\wF�r������M&������9<����$u�B����o
��g7�Wo;��y�{��(�D��o�t��$B��s�:֟���ƋQ@�:�54f�^ˋ���g�����0�d�����WQ+{-�w]V�b�e���k\���?8nr�t*B�+a�������W�����4?�?Ⱥ;���Ǎ�K����_μ/�7��nV��$�<�x�-�z����v�he����[F�>4��:ˑ�	l1�t��W�{8�\f���
��HN��8�����V����s��\��B?�9x���d"���xv�P���g�Z*����_�e���1?(,��[)�b���aWD`�3��U��}@�i�	a1��r��%	�dIǝ���q.���H4H�PF���'j\c��|T;�} �ĽH����M���#6,a�K�W�Z�S�ql=�>�|�V#�"nH����Փ]��^\l;P�qdK9W�:K��lq��dE���mo�M��Wq�rȮs��c��-gt�Pqs
�����n���&�"h�]��E�[s/X.P]&P�6�VU��?)3V}�XC��w���w+��t�e��׸��c�Pt��헞���� ])��YcĝE�X9Sf����K�m�2j��n��⺆?v�6��Ͱu'h�����IX�<	]p��=#IB�DOWW��W�66���^�S��p�r��2 %P�z>W�'�K3����})Ar.n�}J��]��,M���.��Yc����}Բ�� 2��)�{^��Ό�����&��ഡ<YͲ�Q����Դ"	�6�6��rǥ߳�1������3A����ˁ_҃�h^i��sJ�t/�^T{��E
;�������j�����~�����P=�� �W
�vZ�[�}����$Cm�E�[ş�é</��/�y���(�3�L����mU
"�<$��� ��R�}AxڱPB��=���zQ�#�^r��
*��诤�=BS_��-�7?[�������jܣ�Yj^J������<�"'se����ف*��x�����T|	"���~���`j�j޵��x��W�pjB2M%vy�wb���Q�v=%HMJgW]9xPz�����2��U��������?p֢v���?���9��S�-=�¥�~@e�z�Κ`��WL]��-~��� ��c�������CLl�ө�
ɁG�-��Or�,j���	N �>�����p)����c�-N �VVVY[dD�L��}���r&XI��R*�"��Q�J��=1.KΛ1����:�TFs'"��O��Gy��5�$��
��vD�P�$�[��1���p��ݫA���bl��t�����t�2boΡE'b�!�䄈�~����e/�1>�	Y���$5A�����3��[[[�h����ZG|�Rc㋎I��ӻ��w�Ql	�]�8=|e'
!�'��qK_ER��|�n� �]a�"��`f/��A�3�OS�����M���H'�����2���a=�_.'�9BqL�&�������ߟ��2��=L��C�z6H�q'�B� ^�A�ޠ�cݤ ���_�ZQF}x�~3(��E#|�B:�yD�{g�$� �к�y�Z�# ����@����a{������k9T^ޛ'ˌECY9�V�qr�uߑ�P�a��¾�w0�1X��`�oM(�W�V�@�N%~�����P8J��꣧����/v4��pΘ��~�r۠�h���|hh��k��}�o5CX�ÿ�;J��'4�G��0G<5;�i�ÒR�8&|�I�7��\F>v��`�l��V�M^���P
���S(j�/�B�Y�6��G��e������Y�ȇ�6Mj~��wP����3Q��T��$qH�h�<@b0�wǤ���=�߼����v5��;�W�W+��M��Y����{-��>�V�*rV;eo�톇� �V0�>�
 � /+w�"ؼ����
�^�k��s��ǵ�9�9
��}��Ts�j��
ť���uH =��/�vD�gǡ�f�=�O�8����Tm��Ν�t�V�P��Kܭ�!� �5�� �oY�E.��Ì�$������y`K���5*�B$~�.�ePz9����mʟ<ol���W�kFմ�߳��>fd�3xb������gM쬻�j�AWkkk�j�}� ��&Y����\�xWM9њ�?�`�	�$l�cnză}���>SM�c�P2bPeSd� Ҽ4�MQr"X��]�2}����y|OY�\���!����@D	����aP/���O���1��손
Aj�-�U������F�n��h˜��3�1.���A������߽�������"ɱw�����>#�R�w��Gv�Tn?��]T{N���a��J��&U�]�����i�L��?(j�@��)5�hqZH=��ߣ;2��'�h�2�R?�s��>���Uȫ���sŇ�>�wMw^�nr�3?�g�E	xez�t����"���%�i;�7�Z�%��+	�~�;35� �}~��lOVb�>�.��&<�����H�Z%�/�T���|��S����o��#7��x�#�Ub������'���4�R�Idm�9���K]�~}�e-Z�KC��Y���ǇQ\v@��8�5��G���?.���ߐ%��\���eQ��k`�QoO��ء� �� �@��^��Ji?�τ=T�Ɏ�o�@VҼ�F\�a���t��Z|�W)C�h�:¨*uyf
�<==�E*-l|pb�Rv����L���E[~?Q�=��HL�5P�	r	��s�|��Bl��鵐���dOi����e�*D=�Uo�N�8���aq� �x�䒸=�M�A��ǥX�*��i��~GP�_I!�"=�/�a���}(�����z΂G�����A�۪�ǝ�������`�}��=oٮ�tR�r$�8��}*l{�S@_(I��-�M����$Y�b8C��F!��fz��fT�W����BK���&�����a�t�y뇜ZX�����.�������B��,&םa�d�wƓ��<�	�����CJ�����@4uo�s���13��uo+3e�pPM�Q{��E�i;o�l��|���C����u�p�j`dկ�`]����(�Ʀ��ƴ۳�⣣���ofgg7eګH�i�K���mo���%��#sw�`���uf:c��pYR��v�Q���i䦪T��c��PZ�W%���-�$��`p>������xk�Zu�By��^q��?�ŵt�K�@��.��s�悙Y��d��ʜ��1a�E;}�eM.i����cIta��&���1K{3�i�+��z��Y����ڭv�7��_hGT�J*�k���p�?�G� ��]R��*p��M�攛����6�SE�jŚ���P�������9�z�D+맭��H�-��� z���*^����Xt�8��C���M�6�e�U��XJ���rQX�%��\�2�"� v8Tr�|�b�\Ũ����ƻ<�亶1���������'ȭZ[������R�7-��w��WTRʐ�F�r���-��ݸ&�`�o�*�������/�o��e�c�C��M��efJ�Í�2[7��w�jD��m�kBWv*߆��<Fޗ�U�m���<1���O�.��U?2M�����4�"gZo�����a��n�G�6�,�''���(�{�r�x�F��ɳ��0�;�(=CFDP���o^
f�E\��m�#��1ր-��z:|�hՅ��8d]XD�p���z~�<D���p3��|����6��/՟�B?�u����loo��2ˠx4.;.�WQ;g'�9�
�{9,�&	�����ʣ2�-���iW*���~�*S˩@N2��%�)O\�������H��m޹؃bE^^�F��b�+=�)$�:���1��=��f��č��r�׸���O�oD�A �Fj�?U1�)6:�\["a������� f����p�\v빨��4q		�����U	�i�8���Cla�v��k���ME�����e��}��|� 08t���C�uw����L�o#� [���/��|���w�M.檒�����e��)	ͤU��wԴV7�sB��d�!��!�6�)�����e�*i��[��(���;��u~Y��kPȉĹ���X����ICkŀ��x�|9���� ��`��N�2���yv�r��;�|�M�k����b(��4��K~�����Ԉ}�\��J#}o@�k>�LS���\A�f���*��k.WeB�-������PE-e�6"��J���W�ª,I�#֪-O�����(�Yq(%O�?���Ҋ���/�@���#�!���G�ePr�9�xK�d=�ѽ63���G��-+�q����'�Q�O�&x^�(�w{6#���!|ף��vN�̀G��!�A�T�1P�"d+�p$�;<�=�U��9��C��Yn�*�{,I�-���x-�o-�J��.�H����TF�dt�'㉴�\�Y�5_O�#̺D�T޷˹����;/H���-�\���x��?Lc��x�`ח�2�_W�g&�
�zz^_����=� �#�|�$}��ཌྷ��]�=�Te[-+j�V���2�KG YD��O1t�^N�$d���	��z5�"J�p�q�H��
��_ *V}���m����H�Zzxy���[�i��sU���_�����o;��%͵�M�Lu{�M.s����@F�ޏ�y�֭,))qӆ0DV���2*��|�����>_�e	R"p������!٩�^�ՙ��J|�⳽s���s����Ã{��7��`��ڙ��=�n\�N- ȍĠwRbxe�+g�9U3��;� ����X��O��t5v`�9��IL���]Ff1$���w��*��Un����i���㲰�N���x׷;6f�?���DM�m!��HU:�z��$r&�gf:[��h�����rI��p�U�F��)�@��,P��(w�`@"�+���ᬛ�d$ �o���CW�����|.���]���i��a�l�o/5��C�.�ydb]��ǭl�a�Ѯ���f��ٛ��N�a:�����uOlVB� ��+��;J	��DGsӔ����(e2�\�A![�T��XY���>0V���;��;ލo�[��sqgs$��F(%�	n^"���hC[,u��y�l����л%�D�8��򘭭Ɔ]8��جm���"2X�pl@��*�L��Cb�7t�)M.�1I��޹�;��湴(tw��{� O����G�bظ�����5/v��-�E�o�-��< J��'�i�a�����s���dBsD���[G���0jj�93 �/�I𮄢�ˊ\�ؼ�p��a hW{6a>�HJ	��a>�!Q�hƬE9�=��J�E��9�UX��_�2�ѧyİ�����?��%r%�tHA{4^�hO���$�q��`�`�O��ڃ1^��oa�		�6.ӳ��r8���2�9����tC�M85 �r$�!Z�y��|*r�������`�������K��%XO�����ə�x�_?�u-���W���垺NK��P�(T�PW�����d�X�����ͧ&��Ue����}����9�q�V�	��:�?�	�1�vdjO" j�}+&uyE9�A��7��X�րM뽽(8��yu\��n���**%HS=����ϯ�_4��3�.�>L.m��L!jx���%&,��0_g�Ӂ�ý̺q2x�ؐB'��g��x-1�@�tn�9�{���:3�֞ģ�*AX�8$<�J���C��]OH ev��p��ߟ=��88FpȌE�K�����8�+�A����\fy�*�25��CB�{�`�֜Ƚ`k��h���ڠ�>F.��X��Ǖ�[�/U�V�#��\5���yrFV�c�	��ԛ�Er�k�'�f�jyg2�\Ja�;���;���LF������k�D��gڤ)=I�+�$#&Y4�\��2,�"������y}��/V_���e��A�=F�J�բ�b���tw�中�(���T��Z����uO��&B�@�����k_���S{|�RE:Ƚ8�vPԊ�-R����}ɪB��������̪�X|,�uR �M�@���ܾ�� }X�<2�����/;뛫��ڎL.z�
�`��,1�~}&9�j	.��B}�D����n2�Ęa>s�*����3�f�Q0�02���ޮ{���2F������IFN�Շ!����I��B.���_���~b���im��Ԕ�����Q����K��M��1�'���ܰ�<�좝��e��xP(197�kV���1A櫉����]��f+g�WEFR}/�"�Ϣ\�_��>>沕4�_���>3��*�M����VLX��(�n�0�&�,eR
�Il�����|c�bӫ�.�9{� ��6�1���޽�M�UVݤi�p�����"��&��g�m�m��ZvWI���]f��R;<F7�u�cG	���N)���DP{���,�;Q�1ŵ*3,Y{�EZg�3���x6>�p����I�B�q��C�������_x{ �aW`78ڰˤm�װF:Y6�˧����"��Q6r̓��+�/?��7*A�Z�!eOY&����t8v��ƣ?#~�ط��	w_�dn+/�R��%����̯�ԕ:���+׈{�R	��͵�s��u�3|�P٥K֯GO��c�_��F8k���_Snll�**y�d�86R{����� e���F!��u|Ճ���*�_���L����=!�P��<�M
♥Ƒ�v_O�!�z�Nؘm��Z�:��������3��J��`�"_e�
xA��Ӄڱk]ZB�ax��CZ6o=Z6����'
ꥧP�\n��Z'!�:r�C�����8.=���o��yE��I)�o��A�K�D�2�K��#ĺ�{���K���u��O�y�P��!�I{����7��h�HXj;�
�D"q`a��Ч{��DP�\�ȁޗ��� z������x��:����8P*
��ɐ�����h/��M�{��r����RN���T��x�oM�H�n��"fE���UY��ŉf�Z��zRnq�)5m��.�	�F�P��U)))]ql����`h7i-%��S����$U*�m
H�/�6S�{�%�?'A��*�C�U-N���P��˲%�?'��-�?ꬔ��i�����J⮉{3�a<�b{��?��Ѳ��iEh�h�.Q�Z���t�%��J#�Own�1ne�����o�h^i1-	UlK�21�Rq`��r������dK�π�C@+͚Q@+�N��t*�1 �����րɥ6n���n�qG���9G���"�Lz,�:<���`�b8�f�dH��P�&�Нh`�gUr�g�����ͷP��A
���]�r��}�[h��� �0e$ɉ{yy����1�J<�E�'(K�_���9*�y�1@mr�p&���S)i6���mz-�V��>��3��!W�RQ��]� ��M��~����E��2�e��0���ѿϟKb8q���R�~����ǻ3�sp�j����:���@2Gw��	���n��4[����~t����/*�Z�X�l����l"��}eڽ�o&絼4":ylOMCcȭm��$!�>����G.��\��O��zﺓ�>�	�AHL&��YZ ˼;뿷����v�FL�1a�%҆����Fi���W����g��3��v�o'\u��8���L�R���Xg�񭘎c.���K�0 ��*�����U��w����\��n�07ȷ��5p��E��m������-��,W�?JB�R{�@x��S�Ϯ!�q�'�p�ͣ��/EJ/0������O��:VC�	�B�zWZT��!��s�ƵԬ&F�j�㼑�H(Z,+(֕�<6�f�5
J�M'J���������YX�W�|��炿r���9�IM�Ķ!�"�%#�'HDO4)�M�s�ZI�\�w�%j��Aj�V������QQ�M>OP=B���Q�H	��S+�X 6���{;�3�|��=�Ⱦ�L�)�Y"�ʨ{Vo����yT��5�8of�~�]@����m��>_��������ꠀ��HM8I��Q��{烳���L�
2Q�PJ��"`L�H�� ��\�^����T2���1c�&k�t��unp�[тH�Y2C�ED��� Vь��L�ۦ�nY�D�����ӣ��Ǯ�7�\����~ʐN.6��VMy���9�<�3�-Ty�t�����'�FUڨ��3�֎R���3��b�.��{�b̚!QJ�2�?�:p�2±�;��Cj��-��sc^5\<ff>��ͩ�Ð�<B(8ē���P��j�'�ʚ���ر�S��xsZ%C)��HqoE�gʃZB����pq���L���qե�4�}�J1��xG��Ho;�=�g%��L𒷌\IBT�J��Xv-ZK��
A(5o���?�Z���?�d@8�����������/9���Q̏3�[�0qFU���i��G�4X�V�k����1����_��Ĝ61x	"��ॏ2�S���;�D���K�L�
����2�썣`/w��a��uŞt����I��o*�s���������&R�7�Q�p���g�c�ZM����7:j.��������y���#���=|�T���ln�00�l->+�|��YCeN[�=���*���Í��I�����	g�6dQ.���:oY�רK��|�e|�L{$���at�?��[~��R⍞Q�⒃T⼨Ó���l>��R��S�si�����&��y��r���s`�x-=�'�r'��Zl���}F��ٱZM���Q�C��/�zKb�ߜ1Ѩ��֟�����۫C�5<��/�����֓o��V Ӡs�ٯ�o~?���b� ��(������V5D���ԍ�.Z�מּ�|�)��[�K��y��f��ɾ�����y���yK�]=��ɧWxu"%fb��l��IH�L�|&�^{x��ϧ�o��:؎_�3fb2F�3�y�'H�v�<l4�������F��wϯ�a��tno��f�6���ϮJb���_�����Um�Y]�+��<Gc3V�L��������Ɔ�d���"��w�=�n}̻�ˆBN��/Ǟ�f39�O=Ҡ[��лe���a����+ꀮ�[哺�Na��L�c�eR�Ѓi7W��[��Q�j����5��.���a� EW�\F��s�Lv*�ҢFF�Ӧ��Z"xW"z��Ը���a8TZ��O:W�ow<X`v9q�fs����:���J��
i��h����-#�;.Ksä-�em�9���ȕ��6�ԁ�*$d>�S��oh�������]�Y��J�M$T��M-V�N��0��|--1���gZo|��g��=]�8��M��4O'�7���+�=�Tb�[A	���^h�L63��f�B�"SM6��Mh@��Li[zEUa"��l�j�Rz��>	;���yl�ړ���%+�*�-m�L��N��ʰ�𘎶��j�7Za�߱bǛ{��U�CJ:遲&+S����09�&�0�A�e�*���_���3�
L���u��d#��d�WIQm�lZڞy{dRX����2�{�x��M~��ƚ6`��zs⠏����OlR�����n��2���L������)���ɴ�'�7���U;��r��r9�OPY��Q=�m�_;�M���t-p���ڎ����g	CrR�gx*���>m�_��Vm��w�=X����&�g+����q}��b��g�+T���GO$�+L��J�������O`f�O�~;��9O�<�PIP��@�>�����H�����u�X�3_�%���j'�YԘ
K~���,n'�׺~�.=u���k�	r)�9d���˞��CG���?=��������(�jy�/���ϖ^�Ծ:�![;��w������O��i�_��U<�r�'�Sɛ��Y����/dB�J��k'��Kk�e.T1��p!nu�y�_q�����A�YW߄� r%�M<���N
��A}{n���>廤��,�0�e��Q==�-K�|�8-h��24[Y�?���99yp��J��#�t<�Z r�
��L%�������r3B	4���.l�\���޳����	���2Bsn����S��9�A�(���v��<�H�o�W�/�o`n*Z�>�P?�������/�P�� qm�Ζ��� �xZ ���<��K��c5����+�/� D��^���9����;��m`�v[�}~b�p�=cT馁Ř�I����m�� � B1�°���N;�-�ϯ� ��%忋���.��7't��s�
gD�w��
���������\�,�����9�@����^pD�qڕ�W%.����B�tP����RT!Q�/��;�T��?5��/>��D�5��r@�����#~��뎾 j�!_\�z�>n=��V��  �'g-%�r�d0f�BOA@l��	e�Ck�ʑT���W��P�# >�Y:÷�:�Nd��)���'"�Ků�W��B��dea.�XPe�Kh�o@6�oZ��ڗ�;�1��Zj�;T�+r�R��C�0aή�@��@4�ffg=Pb-�~0�3Ǜ�L�����2���Û>�a�,��b�l�[K�x�p��)���J����<��oʺ�
'�\v�
n� n��99x2���,��k]Ӡ
�c�p'��*}�SC�P�i�_Y���G����L�d�Q�eW�!I�iH�-�S�'}�/7����s!WzG���z�Ç��|��LT)P�@c�塧"�����ڲ�j��3��v���TNC?\��z$�Uʹ�16���A��~6�C���z��_ͽ���������^�H��L�}�P��*y ��糆MP��_�i�P6x��B����d�?���B<�XDT�DL��VYb���u+?�|���%s
�H=v"���Z��M�@�]��(f��3'w��F��1��s�J�����8!2š��X���~T 4����o��}�{�����NE���RTg��u�t#R�k�@��PA�>�:�&:�#p����{��  �%�e�B����r@�<��{f��v���R�]�~3"@a }�h������=c�4�y��u��񑑑^��!��N(�s��Lo\�=v��fHd�^��_�\���������ݚѽT:)��A�B��\���؝JJM>�32~��cg�88̷���a4
j
p�Vf�R��L_�$m5�iZ&H� ?>=+
g-$X^���X�t)��pi�2�tqؓ���5E�XS��'��d����������+o�<.�ZR�]<������U=X;ֈo�jXn;��`���M�Z��Qdj���%�)8�֪����[��.kH�A���c �j"u���o�T/5jYyG�V�Z>"�����{�vS��#ކ��:߸z@�H�����̭��¢Y>� ����~���B���\���Du����/�d� �hsTy�#T�ݥ}')## Vb�ju�"�tf����UHuFA(s�$�"bs<���و�Ԩ���5�#4�P��T���0�I�Es�tOnD{���_�H$���R|J��S����cZfZ��2<��[%Ƶ��n	SO{��Qi�$�R�O_AH��@��*�˱���b�uY�KF� ��e��ūW����2��E��*�����X�t�&���v76��ӆKļ4cA�|���5�UU ��1/S��̻�`��#Ź	��5$�"אI�SThI�%�}��/CQVUd�VN�=KՓ|�>\0��z�������O�.J�d3��W垾r������N���{p���Z�`��]���q�P&�(�2Kxa�� �z�*��'�>6ukҕ�.�6�Ǚ2sT��
��b�#S�.��(iv������i� z��+��A~��]Ç���|嚥Ç��+)��O��T�8v���`�����ŉ��`�b�x�H���߂,Nt�O��X�FFF�sJ�c.T���6Z6&0�5�"`X��7�<̵��*�,��"|+CMѣ����i6a*>g�e��� �#��|o�ẁkݿ������?�5���Z�W /;�.'��S�s����}x��"�U!�y��צ<s�c�[�������ڕ����w�y�p��w⤔��Q;4��E`DV}�\�µ��O�L�I��6���C!濌���>����[1�C��|��/��/\#�u��1D_�cKZ�I���.��.���@��)�=' uYy�j��b�1<��K��ݫ���SS���
D� ���>Q��P_��*5W��,��d��H'{��Q9E��U|��n�)�ѳh�;NB�������I�^�wƟ�R��<�c���p�V�HΫ}0̧Y�8��]mW����j3��)E�P�/}� ��¢j}z
�g	i]ҴY`-����>��+?��[����ӈ�e��ȵ�2�o��c�pD8�~EO��u������>"v���Q��|�8�#j�����K,���7"�"�>C��0�,���8I|(��'�6Z����+2� �mF�����`=<<�_Ƕ���me��^iQq+��P��E��y���Q}M\Dg�Τs/*kwA���!�h��_b����p~�!|�7J�?&;<:�FU��-��m�	�Cŉv�c-��p�rB�9���i���!)n�8$�/R�s�i�5+�@L������%u-1o+��z�!Q�h>�����"?���Y٫FT��F��n�q��|`�=�v���;�<v�S��$�
QUf��L��9����0Xje�"z����~L�0�\��m⯵�'T�	D@���O%���� ���� L3Hg'd��2�7)�Ϣ5A1�ث�x
�)���&e�x���ƹ��.+g�X8�F�i��a}-�4� B#[�Ԇ=���*�������"��-ֳ^5]ڽ��$k�Lsf����3��z��h>�3��
S��do��NW�����̗�����ʤgd`_�χ��F��"�PF�����h��c�b�$4��3���	t�S��  Q	A����#��p��� ?���������DךpUW�_:l�q�[���ì����c��2�S��A/�! �䈉t��F띛':(k1qO��ߵ�sy� �PT�^Em������{��	�cn�4�%n<�Iz{߽_�B�"����o����߼O�o
�;��\+�V?�H#Tv���?)��v��II�T�T��lI��B5fj��w&"�CV�v�=e
&�}0.#�ibV�X�Êwc�CI&�s���g#ͶE\�Ϸ��,��i7\"�I܍���d��v�ԯ���K��Y�7ߓɆK��nP�e3���9�a����%��O�4dˈI�}�p1�i���ͣ��׷K2P��Zn�z����\G7�����ϯd(G�OduJݽG`�1�o�k��)��x�����3�)�E�:��_އ����LGGFv�f�����&ǃ�^�pz���W�j���@V3YI��*��S�#�x���Kk2fX��%Y���&/o�#����|�����,,,�N�bHo�FT�g|�LO����Z�-��T2�	:y���"�o�l�|k^vvv�of�1�п����(���I��0ft�ԕ���O�b� [��VL�;\�O<[p.,y�S��"O�x'��$Ðz�:�a��ά�|��̞�D^Q"������&�gb�D���>��z�@%��;��}DPh�Κ����N)1W���6�?�q��PE�����K�|��L�Dcz7�E�B������Я���t��k��9�JO~!���.%�6���I7m�\e� �Jm=�P�����Fhfa��o� gTF#�~����'�sȄ6���5g�1`z~%��A90��n�|��}���3��ƫ�?�wށ������N���_DZ�o?F� #����;�^�-�����;W���'q�v��$��YPI��L&�7Y�Z��!nf=�@�q�"�o��yH��E���\m��:�ǧ0���?��$<�[����ӱt��o��y%{R\�`�&d�ɂ��ړF�[�1��͐�R�~ɰa���E�/�Hk�'R�ȝ.�CnFl�XXX(�0D6l/�v��='Ҵ�N��Gb��/�PvX�	<���Br�T�y�����w\C��[ù?�	�N`��Na\N��Dʐ>�}�IeÂ>@p���#������dO���6��s!���NrI���7���&*͕c��H{nk��2�,�K ?���7�������������D5(���W�����~���F7�g�1��6��n���n�dw��a�� �ܾ��y���mū��
�>|*~"���1{�H�7����*�	X��a��x��I�����7��,�n!g^�X�Ί��4^���$;�4.v��!����[/�F��f�8@ʒə)�������j�v���D�ؒ�?������6����wk6�h|��c\��(���W>N�RQ[Ƚl����lkx�O¿�Q52zw�{��{zn�I&�W�V|���l3H����,k~�#t��;�����������ʝ³���<��@�K�L�,���]��F��9�\Wx+Z2�� ��;�����.��ܔ�|��Wzv7����_11��H�pQ�������b�g�����P5�+��Ǽ4����?s||)R�Db�����Z`�};��^2��8�����[rx|)bGa�9�x� ���Ͼe��9��9О��Kq�=L��kpȮ�:r��F��C;1�qv�"�rx|)bS�L�,++k��0(��)λ�~3���5�����������EDDDDDD�J�""""""""#���`��j�~*���7���(R�N��wgo��P����:C\�w��� b>N-0��S	L ������3ϓ]���S��@�q�Ì�e�ǩ�_��(�HԚ�G�Zw��~/'�n/|.�����@��w��}}}�������%H�j�ҩ0˳��W�=�~�pq�{�W����m���������Ep6��!��1���a�Ù�1c:�$��M ƾ�+o�]��1��i�9�q8�hZ}.E�Puu�h`n��ܽ&����^����	���.�?t-���QH&���7l��������_��-�Zt�#    IEND�B`�PK   �e�X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   �l�X���k�� �� /   images/c6c89cf8-e908-43a9-a5fd-b5d85c65d9c6.png<[T��^J��C�U��;$������X:�	��))��.)�o����3��̻7��<����(��B���ee$ރ@p� �%����1|�����'H�����;ux��IR�I�����������deg���������"�X���J���e.�'�Y�3?�C.;�_
�UL�-�.�Dn�;P����W��MvhvQ����	Xw��l
"�B�F�67�8T�H�U�%Ϟ�=lg�\ޙp~��j)*)��x�x�3�w١��x���;[�	TLE���B��w(L���=aq���;�̐�T&@�+ŗ�V� �X� �7��<�8$��#G��rL��F��"ޠ�3g#3w��@��Ϙᅪ ��w�>��]��_8a��z�=��yffH�I4��b��O���U1�]B|(��H���΢��,^쿇�{���_�m�A����X�L!o+lj�<<�HIML�+��*t�s�|��Գ�M((,��������Kan>�G�PX{�ߋ��+���H5eV��l O�d�����I�"�S ��*���E|stns�������W�ۅ�G~�]di��*/�B�̲�������Mb���X٥��[�Q���-�����!e���֬�w��E.�Rz~���ɴ��i[-����k����x�	�^:���*������y,\��^�.�fߠ�|qҌhҸ��k�ă/���Zb��>���+��5΅2��M�����u^��A�1����4���հ�dڲ7��}'9t�Ɖ�Ͷ�s�Fg@Q��r��e �F�q�U�ՙr��X�O�������uN'������-��X�U���ڠ��:�m	
��v��U%�Л��8餄�^N��PK� #�T�Eq�H�����Zby,�{J��G�����T#��Ѕ�{%����jS~��:d�o����Cu�hM����/FB73�߻�a����Bd���t��g��M���:�=�m��Û|Z��=-���T�����)��󿅘���l���uHS�$R
E����5���R�>N����ʹҋ��{��C�ʇ�/a�ޘ�{��aD.}��ݥ�̇c�� d�~7-(�93����t��[�����&%�cA�?C�#'�&?ޏcWr��-������R7�4�J�@n�ݔ��ߔY��p��$��d���i���ߓ�)�	}��
&sM��"�6�;B��gE���q��/��t	�;@�7x�-� �J������u�G:%�r�v�ke�ץ��ΆZ�_y������>Z����F*��Z�HúvcY^�n$���Ñ
�{��jw^���p �&s���X�?����w�@�[�<�~�`'�s��Y�ނFM�?���P�L=_����Y��>Ⱦ��a��H���4��v>�Z8�n��֣��O�����#�e��L�qĿ�+�Y�����B#1^�.�j��F�y�|;��)2)qm���&)���׭��ND����J��8�M�1s�JVk:��fO�2v�!����RJ������l��&y�h��W���i4.l��eq|�s$u'-�'?���b���<wA�1M��e�������o?B���Y9i�U'"w��`tQ�9@�ٚ0�M5Bs�s���]�0Z������=��i ����g���шo�~�
{z\������55��	 g�&p�@ZIq
t�H�k�w��7,A<62m�%o�NAυ����F����x�Fj��mW�JB0�l�o�?o#E'*�A�z2pq�!%-�����S�W!�hrx�AH�o�V�\�0���tI��'���Ϝ�fb�Ri(����VKvQQ���rTt4Ɵ�v�wV�+�*�����ZG��-�cF]�x)uZAT���UZz�����\t�C0pN�ILr~�Ɨ�>=ea2��ʢ�M�	� ����<u#�\��L�{������sv��B8��+&A�N����5��K���F��~o���ȧ3� L˅��� L�;济��٬@Xorn.,�ߵg��r�0��'�XoB}�T@��@r'���Z�b��כ�5Q���B�M!J[��"��[O� ��Y�	�����U����
	E[r�X�}���[##	0qӼ��W���O�����. ::��{�,���Gͧ�le㕵���ҹDU�"cb�!�$	���"_��
^+��|�Ĺ�����4�Wz����8���l(�լc��\���J��`�1�qS�
�>H��/�ř���R>��e�j/�p-��d��Z`���Vx������9=mdj
'#1�h��?hoj����41��1AXTlg�<��{#���d�G}�5r���ߎjjj���"�bpȍ�c�0<RRN����+~�T��+u�DJ/,3�41��F���0	������ʦ���ZR+��_�5�ׂ��G�����=����H�v��#[�֊S?�^XkW����x����֖��봻�CĔm}�;��rF��������D}Zj�v-}��#�	��i�f�C�QH}x�am�އ]N^��०��іz�P�8	�;�Ѣ��/�%ϓ�����z|DL���1�w�:�7V�v�j����kL���V��D����<��S���Gl��H�A����Jbs\�m��SU�?n��%Yi����H�Nu��:+9���J�Q�vR$���L�N��"���xb�q���j� ��n2�I��b��J0�}:pc�N�㟘u���$Z�����Fk�76�Ң0v�׭���p����r�����OX{o��� ��l	��ׁ�
Z�.6�|��Ƥ���}�l��n/��i���q�I��o��ع&�Ǐ�z��eI#�=��+�Y�R���С����u�u�w����A�ق��|�Ր��~��'-�k��ϟ��͓v���2H��^�Y�b�>�!>�,^V4�O�%�d�R�ռ��u�YCQ���{9����>�D&�8^��Q!��*�-9���mkOOO[�����W��n>0�L;9��Z0�������ҁ�Ӕ�K,$�N0�'6_^�Y��ɦ��ѱ��l�S�� �n�@���&z׊���n��� ]�O�p��(�`$7Q���D�v��D�n	���*�;��zk�%>�W?�=' t��65	��.Ӥ˂���L(����ל�8���_�z%Ze'�c�')ՊEP0�R69=288OH�1��X��	 ���rrr�%s�QPP������$u��]^N�j���!kr]vlddd�y'�5}t�t B'������/��r**�vY�����>|zZ5I͐�����nPD{������mu9
X��m�{�E�٘/��D�E��0����+RNNNjaa�s�K��g�َ !_\�k݁��睙���.��iJ�Ɯ=�(�X�IA�L{��洟]�	����~8ڂ�Ư����n��S^���YU�UY
��N~`g�\�t_ߞ�lJ��BJh�'~~qo�ؒ��2!�d x��V���zJ����y%�tfi�&��7�Qz���X�fۄ笙�������� Ck�D4�<�s� �7-�Lq�������k�>o̕>91������[ݸ�Jٙǔ��舍Y��w�Z������4w��(7Z�fGP��}�"A�6�����	���G�߭��v�;���a�A$m�b
?	��Tۻ�*���Z�Z2�<��.ʖ��t��-�1��d��0]�l�ǵB֎�S��X]K�����W+O�	�����ϲ�����/��a�Y�`;���l�$�)Ds~ٸz��;�	) �{��.,���i��8���i\\?s��r�W�10H�{`&j�bl����t	�yN���:�#�m$�)t�v��cucZ\�M�Ĉu)�B���3�-�@X�T�l69nC'�b#�oR�mƚ���k�w�j������A�%3��ݚ�&�:�m������㽅��b�%9�s���~����~y�1�7��|�I#.{�j=�OY󭳌.�jY�z�6����/Qf���}��闂��H���]�vҫ���ԡ����@6.��:����/z/8k.a*��9đ}���eЦK�TM��l��z:<�p�V����J����d�������� a��`M�bєGR2�����.�SQ�h�,�3\�������:F<��Ɩ��w�����u)�Y�"#���D3zt.�^/%��Tge���+-��Rx�#��uUT&kT3aa,uv��L��'.�#�I��!I�pX�ʲ??��3+�v����X����@����R7�����Wǫ��~c-(�`<-#o���4���A��lh�I;z�������j�)[��c���(��w��F��&ΐ)����`M۽a�7��(*:,<�����-7V�w'�1b�8���?��c�Χ�9}j��1H�*��cS�G'�N�*�;)b^�HO�ϿM���OkL���4��J���ƞԮwu#:3��㌠�|/�����v�&L�-��r���q��9S@���������=���x���D��F� �F����L8N�"��r�Yf���8;������;����=5����T).i�}�ax���varu�M�(�ۍP��L}/�tdb�gٲb����Ѵz� �ޠZ��V�K
@k;c��>cY�|��s���e�Se��լ��6cbbZ/d��(y&]�h5�(��q~����j!;$$$��'	y�]��?M<Rq�eȖ�77�Rhk��0B4�C9��?Y�$�I8qr]yc��Q�;�����.яT
�P�.t44�=]��s(`��*���t�/[sy@3��W�:�?������f�=<ԝ���Tb'��W	8>ޗk]����r�����K;���$5�����L7�Be�)��u���[[v��0&v�Rf�Uv-Pf:������N��Ij@�-��Xq�3����7��{2�����T�=;�X&?�{x9;@��O��� ������]Gj0��n1����Hf:�9ov�'5��)n���o�e���%�6$GG[�x�E��O2Pw��>�� �.N�����N�T�u���ρ��_ �ܘ�J�_^�WZvx���:�'P��N~UEz�RW^�a�I�\��7�G1�윲���D���s��)]_7ҝ1�QS����!+�����)N(��A&�s��`����ߜ����ӷ��kO%Ɨ�I	l]�M���WaP
��/f��e�X�AU���0Bϖ>��N7)S���h�����u�V�c>G<:�����.A�=�8PR����ʎ�Y^1c��3��&T~m1�5:t�{�F�$�Pgש��3�[vF���U#����B�a���6�e�	P�<L���7����C<�ϧx��F�v?ES
G��]A��i�����d�oO;�k�l��c��a���һw����H:�����z�!�YAu���:'P�ϯ�H~���Ǜ���EN{ q�=��Y���H�_�`�?^��{qu�=����V��o�ޢV ^����RTQn��=�o�t$���@8�������Y�66h���̬�����%��4�z_O�q�wo���,�������qc�8�,�[+�'�Y�Rf����[��'%�`���vO9������éG{��Q���
^�+F(&��T=��.���V�������7�V���BJ����X��XA��b���n�R-X>A.�U!u����+B����Bl_��cGt ;#ȡ�������"���Q^�-pwX���;Q�}EB�7�-�|�_�������v��a��	�;^ב���,  � ��*Rz���?3���a y���N�	d������1{6L��v�ym.����˫4�����f�=���;�}tH��n�kg(��Y�û�����ȇ�U���y
��9|�����Ӈ5�
��哞sH���cW�sʧ��<�VoJ|~'�d#�<�І���&��u��7�ޛ��ݲ\����Z��E�n���H��t��E5�j����Xo�ؘ"���*��rx�Ah����S�����{����h[�a�*o��}	(����zK;;)II����4���Oj��@���(��y��{Է��,Hw�ǗÇ.d<U[gc���_���4�.�&�v����@2�1�i9�A�ǭ�����=��z�0F�E9�xs+�U��AJ�Ί���ǽ1��� Iq Рab���77;;;�߾�����10����c)4�n�W��B7�[�'�S����P�9}��.G� ���[Z�O�[W�gff68>.��#d�E�ݜ]�@ �p��n�{���B�H��z7{5�]���ސ˿ �����͜�'��t�ų�G*H�wt�����/���d���ǁ�l�w�zͰ'�̆��;���"�"��o@0��V��ǈ�΢)��U�ϻ	D[r�t�bf��NN����I�6�W��J�sNz�(�㡅��Dh�5cø��*��x������|?�Ϗ���}�,#�λ1�w����$�jl��3�(,��>��@ૠ �9��� �;�ט�����R�=�Ѥ����}�_Ϙ-��R@�Ꞇ�k�-Y=�F�>M4��'��忀đ?�������ϛ��&� �0�	��C���F�6:"Yi=[�0 �w�X���n�i����<��+ r�����]g��l�UzS��!kS���-����5͗/���^��!��x6"(��း҈`�n��n���>7_4��ܲy��"�g�5��E�q_�*<<ϋ��D�R��B�$��%�2	�z
�U�������ǉ�8r1��|h����5�q���"��Z�����g�9�#9Y�b_4=GF)}��?o��c�w?���!`�D�; U!�fr�F���I�]j�??�r,���w������N��y�u�Ţ����=����-ȅy�wt��_r��ծ�j�<ٚ�� '��}�����҅p�2=�4�Kt�B*�i` �����'s]����I��zt��=��N��+-Ó���6���b�A��y�(p�#�8��VRFL�Ȇ_�Ir�;l��\��O�Ԁ���V��i���v$� ��'M���:$I���oT@�<卌�����O��K��'��d��=��k��㡶�SSa���������|�	�X������G��bX��[x�������O"���/2���st��ħ��F��T�]�!�|zj��⃎b
¿!`V�?��T߲��h˨��@�ʊ�W-��}��g��'������ɦ�<�j0',%q�Bd'3C��}x���h�E��n2�3��7���Z��$e}|yn��V������a���Ub�OGX��{��ou�QF���yUA��7h4R�&D��N�3�+��r�D�M�p��:N������8`�t\2����51��F{��$ �zJ�6�b��B3�(.��9�H�i�rg����;[!��@F*~��&�}�f��Ị�����S���]�������r�'>&��po˴�!�V,�=3��`q)��몽�����{���?���EQ����P��7 ��{w4�58�����Ģe�ޏWnJ�8��UvKHS��K�%ǳt�A�"��5���A θ���*ޢ�T�ۘ'��ic/nԑ��MR-�1r\'���|���{nl��V�F���m�Հp{�g˴�#��X�8W"Up>��K�z�t�BrX��HFmXn�����v�5���&�&m;�g�@k+���ՀT�M��sr��ے�\�`����b���˥/�Z[�FBZ[uN*�^�&?݌O����"{��e'��#��Y�?B�;��Ț|�Z7gt�SF�:�l�ߞ�lV�W��Ґ�w��U�.���������1o9Ō��Jo���!����x>�7���K�6嵊��;��;Y:1�^�5b@UX��$�e���E�lf
B�����_n����z�*?��K���6�Z6��K宐n���,�P��䵫U>��T=P>�4�}��LL��9���Zz{�w?����s;��z�u���W�VN�����~����@�}}k��2\m�\�����ߘڙ�6`�p�w� �yx��]|q��K�L�{t4[!�]��!*r����}5�������Ol���BT��`�'��XZ�h��c�7<���h+��/�;)�o��Ҽ��Ѕ��	��GvR&`u���>�C�V<��|'ח�ll��j�)���'���;�Ĥcz�W�{��E@�SE��B����ws BI�
�0��>Z�y�V54�]X���a��f���7}ďy��*���v�7�z۩}Gif�����B.և,���ln�o����D1��U.�Kw�g[YڥV���D�[d���c�i��e�N���w��"C���W/�d(0� ����䞵u��`���/��?߷�|�� ��Q������7�k��?��=$Oɗ��h��9wt���a�m���R��s��]8��9,�X�������J�Ḟ_=]��H�ߤ.V}��t��_�~��!��4ލ�AJ��GuՇ�\��B�r#��Hg�� 	&�C�7y��G,��:���=�`�A��H���>�{7����sW������g#ɄG+7߸a�pq�\�mJ���n=�(���у��|�$1ޫ�=����{�H.m��e ������-r��qV�����I�t"���p0��IC8��?n�MB�r���Js�V:�)[N:�7�K|��C1�	0�U��j�����;Z�3�����>d����#'׿�zx�kPr	ݳ���%,6y==��h�A�i��# �\���!�ǐ�y��6�<�O��'��T9�5m%��Wr�C3cLs2��<r� �@�z�m���J]-q����゛`�L�O����QBU �+��!R�D4U^~�X��i�˚��tck{���ܖMY�e�"$�����X�7$d��D�RUɨ���1�t��J4':_�%P���R��q��������|[o��{J�{�Rf��-��>�z�24�J�����/���������p��)�|�B��{'[
���b��%�(��H=r����ԇ�4��C�|��"�&�Wb]U��IK��?��deqf�n{�0�B�OBk;�n�%�e��e[�k�Q����z�ĠTR��Ƭ2ֻ�����g�dW�Gz����k�v>'E�Ё�=C��봶*�m^E�rY��?A�X��.y�<�o6,LF<[��c�b�<͡�;�P1�wB��66�V�@ .>�)�y#/
J�k�-�N'K$��<�0�rY
:4��i�cc��`d�g)��C�}�li��P[5I���63�����u��R��� ��~G�+&�ْp����n͢�u�O�Y��SQn����]𙖣l�O���k�^�{�h�+\��̛�PK���:g��\��иq�B�Nl�GG�>�&�
����DƂi��)�3{LqN�>�;��j�)�y��&m�Ȁ1��UM�5z6��ɹ\>��vФї�S���V���u���7���V�	�H�I�W�#��]���ؠ�^#'�/Z,D}7�;���px����B>�Ob�6�|���Z5v��˾pO4f=�t��	�P�
��2�VG��@��FO�$�%u�������D�m9�^�&Zfff��V�r\ڡ],�_.;���\�^���#��V�b-┅�|I���ˤg��|U7��ŵԤ���nn�����J�D��q�!;���<�G�[Hɩ���wݰ������b)2�K|.�/�4�WK�=����䁯h���jT�nTk{��s�(� �����ԍ�����}���cu�Eˢ����Y=���B������b��:%���[���e��N�ނ
�۝5�K͟���*�%����B�ҧ�$DEaJJJ~��SU7\	r�LHKK�mD0o|����7�{KO�����h
Y+J���3�ۀ�zN��@ڒq�|�$���X��c]}}n��V��ſt	#���~f���M�d��z�e���i�8j(*H�}�-	����`Ӣ�Uv� rdÀ��������׊��A%h��Ҽ�UÙ5[�JG-X9@%F��G�G�U(�DI$�[��B�`X0���x������v���
4���/�C�7��}}㇔�oq��kjVNije��P�p?Z,x,�[�� 0&���J-�k��T�Q�yM��P7� K�0S4��uYxZ� ��C_ZZ<�� ����.�$ʖM �F���:^���S�eKj����;v<-I\�&>6�a|���T-���Vˈmш��:��O��x�)��ՖP����A�>x��D�5"|Q��#xV��.��:�-$h�mC���&4l1M�%���~+h���G�B�Wׂ7i����l3���jpLƻ���y�5��a��8[u��ۯ��¾�r�
�@�M�!$��07Jcc�W<z^R�g�4ؔ�C���霘b�5���\0�'����bx�������DPWW�SS�c�xײ�q�#%-=9=,�̔[[���wmF劣`�-��)4/{t˞��� 3\�a��]�p� �z�8biUM+  VI�d�g�A���.�.���<�fZú�T�O�����}�S�(;66ʝ=�Kix�����2i�`�>��~��|�1���o��=@ԓ�:k�c��!�~,$xEis|W� ��A��ɽ��j�nZ����تb$	���/H��ֆƳ�܍�Q��C��fGn�K��wص���C+�~z朴�G�e�k�i�Մ��
��R�� �C��-���y�$8o�x�h�/&%FTek�#�F<��:�A9A�x�'/�{�8�����ŕ�ƽ�E'��n�씆=��_c�O���)�P�Ǯ5H�0ᬬ����v��� ��@$�$ϻ�H���fs�ȾW��l�8��TZ�!xQ��Y)D"ߧ�X����J�V�����/)����ƹ,��j-�b9�}p ���Է�n3sX8bI�eI��������`U�-&8'0%��θ��~�0V͝'�}6�@
"d�-)E�=�a��LO'B6À�nF\PP I�P�X�S5#��Ά1���茲�����5�W����b I	��]��3�¾��+�-�B�Iϣ"�xI�"��PՄ�R� �~����Я1��wh�R#eH='��2>1{�m���4"���,�����0���ѓ�&	��%�?.�e\��k(���R�j�F��(��OT[<	�L;�d=R��<�w)�a����[���&-���ě�ѝ�9�o*�������ས�f����-�������2}�a����m�Kx�-`h�&K�h�]X^�ʊ���}�)[��CבcnUW:�ѕxRKkv�7�5��b1��MZ������<Y����U�xVN���
���P�2�I�~c�.�S!���t���?57a��
f!{нh�E�S�z�{��!9Xv�^�Ă�.SC��A-��|�;c��xP�T��P�904��'���WI�ͣ"��9r�o�濐�V"_�Ʌ��y5�f3l��i	c&
�M��M�6�τ[RZ���&������s-=KJ�]a�����.%���>i:���C��"6Jh\�@���yM��l�����)4����o󣂒R��!�)���`g�e�{::������ki����h�i��.q�&���m�5_��jL���+\^����	����y�� )��;�&�FF��9�a6��Z~1��dI
��R0ĲK&4�}Y> ��2iE�R��y|z��䋃m�8������W;88�J�pu��V�V>y�6�![*+��� F�h��(i���3
!��豰��M�����WH�X���ǎ�U&�N���^ư��D�����]�p�u�z��L��e�p���3�� 9=����Y�>�6�)o��ؽ{X5p�/�F�9��i<��M�����s��"9k0X��"�p��w�*�c��ic��|RG~*����k�tbɃ�(��%���R|����rw��;5M��u��h���"C`Ȃ�w|�ZgxdDYe�_���|';��m�W󓼗� a��O�;���#���)�m	���}ޜ���l�ҹ����B�_	؝xjj�����+�����~%%)}]] ��]���Y��7��x�1V!)Ѷ�Gm:%���%��]��@����uN������2p�0Nx���m��?A@���S�i� ��3��wF_���7���?B�I�i���}�KuG��x|�aI�T4�dX��4\�����P��9M_=�>&^B�Nv��6a�����}IV�ymn[���6�$�P�����JАi��yz����n�k'�I��vOy�a�E���N�09�g#N:��- �ɠ�#<l�۵�N�H<���No��hXR�[�{j�0�l�ˏ��_�W+5�Bͺ�r��r�b����S~�>@�����.2:��C��SwN�=�0��5��0Y��Dۦ�ZY��9�{ ���hɋ�#ɭ,<��"X�Нþ[���֭������߿���-T���f�am0R�=����`����MD?l�b�)j
����}1�/����7\ @�.�����~h��*H8�t@�c~"]�A��}tI	���pk_�١'ð���􉝄��y��T�@Q7��5uݶ�Oۢ)�b,Eڛ��_Z⦖��`bq�s�' ��F�Ϻ���fC��U;�o)~�s%3�C�Ow�M!�����x�n��`ӥ����EAQ1��=W��~����Σ0�����Xqh%!ꮍ�Gs-��w��<<A�
�z�%%@�Ne<����ul(J�[� �������
��H��}�����Ld~���˱�I�<��B�o�]�B��,$<�A�H>u��$E�8��'��v���d&	���T�n�D'���}3����|�\�KK���r�L�߱%�������@J������V���z	�=���,8R����y�N-K�ek ȲY���i��D�W��ˋL���}�~RB��g�-N\���!�qr���	'4
���b���<������_��5��UT�~W����vR����N�u=�{�G<A[�O$�.g�G��Z�4�����������-9b xle�n��g�$xX�`�٨�����̧�Qsq .�W1����D���1���]�"��4ڈ�v�����\���g���|���立�����f���C ���p�j�;�����~S{��F�,|�����߾y,WԔ'����>�9_d���]gH �<3����u��9H�i�\�ǦV��o�)�������sU�<]m����X��	�
JP���v F�r���E��D����ϟx�Ny�r���wE9��}���~i��}�#UWW����)�$`oL��c���J��n	�h*���K��`�cD���UƜ�w�(��,l�:vw��Ї�ה�.6��^V")�R�%��T�?�f̴@���� d������3�PH��м|��tp�ਮ����@��!�{[�U!�+��{~��㶎	�I~k{��K��zu�!��8	�	��j�#�Fқٺ�P5$ ѣ��o�f.���D�T}�0�s�?g�7�\���"�R���4�M7v��gs�oyyy���Z������������=���ЇR�4�[�JM�D
~����y��f����6�C�(Q���G�2NB��N������H�?%p�OOOe�����������dJ�24�p�m��&I-V��`{Ɇ�d�� #����/hr2���T�T�q�������5cJ�MK�K���l>:\: CWӕy����7H�b[}��+'��Y�h�c��{o�J՚T�����ƽ���(�o�egcc�I]2A���b��h�֒9�k���f���6�tG@�j���"�Q!YZZ�X[x�5?x^S�|Drt��杜C�����<����Z;g�MӢ�������b|���6G�y��-���NbR�1 � te���Vz B8 C&s�%y����[��u'�����M= ��p��,�ϛ72���m�|�
��+W�[Ԕ�~0{#���-�5�����];p�W�뽥"�HoA#��� JC�{�����O�&�o�]RE�nd�w���-�l��W�	�1B� o���1����QF��Mf��)�<]���6�~J�ؼܔ�~X��V��?oIog0�¤��g�o5����2�>Z�0���6Iʐ�k���К�
D?`%�Sƽ��*5J�8J`�	�zv E�X�@e��霔��C¢K�/�K�Ȟ?���tp<�v�b��e�Э���bH���u�$�:�>����C���ms�*A��i���#���z�#����:Y,����� ����py*��3T9yK.9--b.�x�Sog�x��"u�0���@0�(A Ԥ�𼰒�����8���j��\�P��ᑹZ�m j�)�Ü�qh�9A�v��vcݮư��ʳ�9_w�v �?���[*�e�n���@J�����i�ĭ?<t�g�
�a�9������m�%UNkǍ��.��+������\7��M�����hx5ڡ�/�X$5RNg'%��>z����Ni:�$���R���ќ�̘%��@		}}
���p��� RI,�Y� �f,�
@$�4��&��K���9�&�2�� �q�G���I�xb��/����������ל-���Gszc����yW��>R�����;~��#��O%:$$�wO��p �����J�}�Հx)�w^�F�%:CV~��XB-%tЌ䊼K�w��s���z�oMF�f��I����||�A�
���|r��
Ŵ��{>�'�ߨp9Y�&Tj��:�kZ�Q��0a�Z$��r�>O�$j�ʇj7����H!�zD;8����a��.9�˶Ǻ��E�4�R�I��5[ު5�t��]��F���Y��^�z1���])��VEo�z���yx�7/)Ӓ���iS�$~-��~|S�bQZz2�[]�Ȓ0��Z����u/!J}ϣz���$X��/YI��V6�v KC���k��͘�i�#�����'g�*�:��,b���@��n�Ն}# ����;=�sp�6e۾ș�&|@iGR�+<a<���)@ũ�Vaz�����,����8��ѐ0��Qg窟Ӣ��X����zxy0~��8��%�GTۻ C�U�B�������L��ܹ��>+)e�T��{s�c�������à7)�.%s�إ��\Pq�H�㣏�wW����6�JO�LL%^���*���o�-�X��Q:���{����쬨d۩".�OŞ��Ԝ0��2�`C�;�[���Z��[]��,��e'�ӹ�7�VC7٫����ٛl����(�/FAO�1?0$�T��e�}6��L #�v&�O-��)��������B�$� e�#)��L|���+㭔��@S��9;chXF��{a��G\W�S7�ۍj�Qqv0|Y��rOo!<?�H߇4�%�����0rtaa�&��E"�鍗�M����P"rK?-U"A7!F���bDHim+�w{��Q�Oz��1�N�$��rBO�[��O��e��|vp/vS�wWj-�������J�,X	"�D��Z�x�!�Nc�D����O�+XT}�� 2G�*/(��ϟwON��$yo���L�Tc�b8�d	l��jȼ�B��a���� �ؐ��I3BNW�o��e�)1%���&����Q;�~6����s���>��G(#�Z���G�l�~�2>, dF�#�8�ITk_�H��Y�����W�J7ܝ�_��JL~��������;��)�� _:l?�azk��|r��Mc�?T�����!��D>��C�/������������/C��Ъ4	�@�7���d�OFe$$��������a�TF��+/)�x֮�ʤ�2@�ot��VUW��T�HJ�*]T��`-���B4����Qr&�����8P��J��U-9o�D�K��'8�Vח>7l
�^{>�vU�؏jǓ^w�T}}�0�{�K��w�0?�yV6�R� �I����.�-)Ot�Q��i{X�	Տ_��C �x���	�=a��+�J���<��o���c�y�UH]��s==b�ёe�Z��KJ��,-!��((��gn,����o*"]r�>�l*�WU��__7H��j�(�r�&T��纗��I���`w���󑓬q9d�"Kt5}5rb2���s^�M�B�����ח1�$xkHVb<K�mD'-<�i�2�����!��a�`�/p���6VVo⇶J���L�v�~���B����TX)�v�	��_Աd��;gx�~�%eT[��J	���b�~���'���bp�'Tԝ�9��[��w�Z���yy�.�>>B
t��w�T#�3��-�.�����)AS{k������~�լ�8N��� *���<�ʡ��&�U��q����U�Q{�����U,>'Kgof�P�k;<��)��mF,B�Ԩ���������^嚪
99�x�/�T��e^��� Y��*��a�))2����˥|�ueh������T�a7PV���W�\(�b]��z��N�PO�����<n�:?��<��n���q���	��/�!�}#U��6�?'''��rpv��"!��nb��e>���aY��i�r��k�c*��8�S�o?��츱����ꍢD4�x�	�����{�ҵ�����ak�NG��S������Q8��0%   �)���%HH�ҝKw�H��t���������+�4�,�[|��?q?���x�2s��\ל3�)�}����p5���g�@���g�u����?9�Suͅ�8p9�9{{1?ʡ	��Ƚ��|7W�l���A��.��14	�8����+T�-�P�#ؙ��xG�"�^ ��������:/�_�>��+&�Պ\X�;�g�����6�eJͦU���1�/���s���8�}+'oC��|%zL 6�>d'�Ŧ�?�7�EYU#�e�p�ns�]S�����!n�S��۬��ՌM1ߴ�<ts-Lw�rt��E�\̠�,e��+;mv�$&)��;��:����*�W�xT�r�=e�zOg`�:�h`�#��8(*��_c��À�g bss��(r���S.5��d;)~D5+��R���U���I�[��&�!���J.p�66=rߤ��nڻsU�>�����wFE�-���J���Yߨ�k4-�8<Oc߮ok���!>���'Y��4m�&Œ���|�%%�\�@G�$�z���N���A������o��-l��o�f"5}��0��������B�H�x^�9
(��w�7���O�{��>���/�+��x/��g�-�`�b*i�7�	G�[h^;�M�#�)Nl1��O���M�6w�0�}����H���n���ƒP:h�.�v�����ش3�Fnv����T�w�g���4�$$��FJ����O��h��%�<<w�.ʍ?��{�Us^Hq�n�&�if�M��QL���'1�L��..�55�J���D��Y���|�|x��d^?�ϟJ0	}lV#�S�Ձ���*�Ƅy[���s��xCd"�@�� ׋���!:���[Dw�����*�/� DuW
��;ks��!��z��b��K}�u:�K���7�y��ԕ�Ka�q�'l[0�5Kc���Ԙ2�6��NJ*�L��m��J`��%�Mlf���wp(xZCz<��hd����A��'�(��gq3"02��Ƅx�6�Q��q�:"~ĳ��%�f<���!]�[tk{�+�4מGw�^�]�t�5h���]%��W�i�50r�H��v2�I�����7��M�k�<��\XRJ��)#��`۾\=��{�4�0�;p����qJv3��W^��T���������& �[�L�������4��/����V�h����k�yR�Ɛ�r��(��c�0�tv����$ͱ+˒a��;�8�r	�-S�kR{��c vՕT�j0���Q�x"�>���Lg06Q1+����%w�70����@�:�|UaW��R`��2u�:j�تΆE���zƞL�CȤ�y\��c�.��Y��B-�9���� Bb)Z��k � �dO���L[���p�XI���d�-yR��$2�w������l
��8̷�&�|��g���Sai�){��&�/����>�
�)�W�p��'ѧN�� 0%�^{��X3��C^�s�飶#ʳ�ǒ�lL�k�#�*+c�>^K�j[�
��Is\It9{�����{�%����dhw��gv~~�,������^4wa��z�
����w'q�UGwv[ۢ ]����%%U�LՂ�H��^��d����M���&O��[�����~���v��$[4y����ag��Y*��1Ϩ�6�Ɋ��̓F��h�)/ޫ$�?gWg;bzؓ��]��ޣ-5Oݦ��#���/"���4B<n$���Xm�`�Q��V?�+(*��4e���Pzߢh>j\2���n��&�+�`oUԯ���v��y�O��I�%�ƶ6��]��m��~}y��R��+�#J|�M��s�$���[��'&<�f7��t�<QSS�1�p��ὀ��k{jj�t������`̇3���݋)���w�܀NȆiD�/'�_��r߿�����n��>'
�vF;Y�%@{o�����z��$y���E�GNEU�Ї鸿�\��9�����Ϩ��`�j���F�0�P�XS�
m�'���IS�4N[��e=y�f���cD�L�ȓwEE��	��{2N���JG����	�h%� C<̿�r�ϟ���W�¢����Z�|�Rz�"��f�-�5	�p{e�����������9϶$=��x��TY�r����$��13��?2/8��.���':0d����S�em㙲E9�<{�?d��ѱ�\b����wk�H�ތ���#>�����NL4��Z�K�ZٺU���<�FB��W�#����L�܅�r�_�D���!�P� �:_��ǖ~ڱYT�b΍�_	[����B���O��Fc�I�����������Vk!�(��+�V����q}���9��f,���FIˆ3��e�GAA������;<[�������*��/���j�7��H"}2�o��<�oY�9��Dz ��\e�vе���?�P%��>L�|�,?��:�#2
����M�~���t$]�$�{t�V�tW[�& �Uǉ{�wX]]MY�_7`�N�Z�g+��#eu���j���ð3���`�lNk/����׹��;g�~����Vڼ������*;��>/ޅ�m����K��Ch/���(W�꛵�ݓ�	��S���&#����j��Q^		����l�%��B�x���dU>�X��kr��� .a�������b�|�����&�[$u��˘��aP����Jc)ë��������֠w&�,�21�j�����ܓ��i/�sB=_x&��0�z����T=��u����t[z::2+ =���is$�=�DC���My�[�'~]*���'��?���K�]����³ؘW����6��ޡ��_$�\�x�#�?������Iu� ����������7�Ȑ�g�-��	�"b߁����I"8��RqiJ��� ��|+��s��s���¾���W\G�Ҷ��a����M�?� ���Df �6��*��`�čI���_�
��ʇ����r�����"~�OH��n*�O	w[�TY�����
��É�p9��@
{4s{��ʄ��
q��W]!y��E�������80��?&�H�S�֘���o��7O�����#j�ՑoE���oc^X��EGs��J�Q�cnC�ښ���B��Fc�]a˾D����k��������T|z�~	$3���<�d�z��ག��W����R*|�U�%ӛ�62�b�I���Ο.Ә���W����9�����]�c⬃:A-���9�!�D�c |}Ih�a4�d��}BG��ǩ7��h,�q^J��O����no�]����%�)e4ėGHJ`ô��"  @�WsT䈄μ<Z��(EGq̈́����"�\���UY�����o��$� �뜋;o�w�o:I��	�<������!���P������e$����ο�u4}C!+�[$�^H�=�u�_  u�$�O��M���:���h�1;��F�J©ú��``����&�dB�P��Jw�/���NҶ .�|�S$��?���OV��=�q¾�
`�uv��+^�����`�>L�L}�f�)&7q�4k ���Wr���Η6x��zh�+�G��R�~�l��&�G�a��Ы�{����u�u��ښ��ʮP�f`GF�����Ϳ��[㜨H���&Y�A뙟�l9ku�DY�.���X;+�\{J[���'��%���7�{�`n!]4Ԭ�Oؤ�{�8�{q�OS6WCMa9վh�Ϩʯ/̰^^���`��IC�9�n���R
.:�}ː�y��Gڎ1c�c���V�(�u}�����9�}��Ƹ�wS�P���Qz{J��(��
�!��eFf���Ò�&�'
������hn7c�c��_��qz�-��X�1�9�4y���㙳���"�7=����Dɚ�=�w��K��`S�MR��i�yp>0��ֳ���/��Z�"����z�G��v3��<�zz�S-��J3e��	���l���mSt�=��d�0Q��K �:����e��W�V"�ߜ.��{*f�N��~b��8����K� L�ቮ�jLX��{�5~�Fwo1KLd�Z�%��`O��o�1z�:Ò�o����=����W�Si���b�7EUU�'���	�="�mB8�O#<�M\��o��������r�m�`��e�8jV��OG�04 4
_�%^����	�Y�s����W�(�h�P#0����u��o�E�s�[����`LGl� ����}���!��E��l���K����WX/ϧ��B&�gg�X;�ӟ��;�^�с����6�dݮ���dx�Z���C���H�	�KmVo!�T#�1]��������_�Ș��`]�R�	&sVyW. ���f1��V�Uf�G-�a=���%r0�jvVϑRt� �i��('����%��@Hn?���xU��;0��W�붅C ����J[B|���D�.��[������~(H+m$?��&((�γ�p�Ǡ��#(hq��IN�)p�;�a���X{}�u<	�տ��D�V{r�%(��ۡ&���Ɣ�g>�A -���C�R�[��s�AQ2v,�PĪק�lڥL}Sԟ@W, g�p�l�{�z�shw��,Wz����-���ڳc��z[�{x��$��G@�!9�o�Ka����>�O��/'��fn�j����[�t��	E��{"�SqQ�W������T���	���0A�W�V�W��1�m��e�o���LLL�|��>��
2�)�|��0-����U_�g���I��ǃ�1dkg���E2k��(��Z���L`ܟt����fڕ+<2|��udD�3R��jQ%[��T�̇�A���Ҍ��6g�6r/�W��j�g��XB��I����n*4��r�8ok=��z�J#^:��t@��k�v�5w�ۄ���}wL�4रr�6#{ܥ�����{xw�04(���QW��gA��U����+s_�%��x<�/�ZC|�ݮq8��Lk��|m�!O��ؔct��Z��j'R�fZ�����N�(r�2�Z�자+�밵���M�55��2r������[B���Vպ��D��#F���r�>֚M9�d1��.�@Y�ۚ�E��FN/����d����]�W��v?���v�` 0��^;�+UcE�ۂ�-~�B�L���I�`Y�HSY�fhhh���M�����ڋ1�[��+�fH��\9����s;9�s��b�k�:������S�Y�L�C���B���E��F���t%��@�&�[��k̋� (��rJ3��Ý��ύ����R�GUF����uo���l��w��b����^�?�(�:�(4�u�Ag�s��#�j��t�I'���Ά��`b eE�2^ѿ@笞Nk_���հdҲ.&��7}���*���"�I(���F�8����\.L|��j���'z�%oS�[昴��ǯG��Ǘ��CV�7<�g?�*���j�mb.Q->>�O�4���	�ﳁ��P�Z��-P*�%W��i�3=�pՔ��1v�~#t��/�c$/�Yq��狄�-5(�M�-.�7aHƆ�r?� �&&��������ܴ��Ru,���/ǋy4&��,�vވ�{s.�1Ҧ����h���k�ž�{����������V������ȳ*�%��:_�B��kPht�%��%D8@�*��uх6��#�8�V�0�`�oΰ͈�W�7>�t�6���)�I��K�o��)��w����Y@P����o+++�62���$��M��#�K g��*�C�s�Ɖ�;m|[ķ9΋Y����3P�ԁ0ihJ7���P��H*�!W*$����ռQ'��\���9,�Ò6���o}��@mF�>ZR�k��p����:k��!&Ih�����+O��o��L����{K��{R�6n>�T]��9gvC������J^2F�>¡J$Qf��@G����<]�����2:�@Dѱ2��~3�����R���x�]��)J��WL9�����8�-�x�'�-�S"(�������ga��#u��XY�Ӛ���}$.�C,��2���2�"�/ӗ-�(m`�j詮@��(B�k�5��-�+��1H�O��n�&��M��d��$�/��FFZ�������we� ���}�����H�3�l�GG?��7�r�~ԙ���!��_]���Μ�w-�����2������-7�${�6V~�آ:�>�,�2� �ikD3�9�q	��b��Y����~M�%�Z��:�o�	�{�qІ�q����G@�r�  <:�=�mC�7*m���[��^Tc�tl��o�i2���+�����hڷI���Vh�{��a�+=�Q�9־0u66�:���tn��S��W�؄8����uy��A�띳����J�3n���.�ϝ����
���hO>�Q�1!-,6|���Lc)no�Z[{��g�4dkY�� I鑙bre��8v��9E�D��K�׎�}QdA�����}��Lq1�G��R��E��Ͽ��rY:�>�k��	|�5"My��mє)ݏ\s�_��>����q��֊d?���#�	�\� ˏjً��-��%�\8�l/���F'FI��}�X�g���.,'Z�#��WHHo>�v_l���9�����|pʸ�������evěuq�����V�l:���U��B͒�/��o3�jA������ a��9��cYMG��������'C�ú�i!ߵ�ѝrd>'������X��_z���[�>�ic�+o�[߂�ɦ�(;���L�{�39^��>2��Бg H���鞭��6+���Z�2p,� �cRn�t�?/��oA�l�#��}k�"bZ�	ts�;ɏT� ��b�<�]w�gTh��T��UU�6�*H`AzG ����,[������_��*[��`ö��>l�!	�q�'�SǄx�^@Gʄ�6���~mb�7��{��.2{��^knW����l�k���ź(���B5�S!��H�?00F叭t��-�gzM�bX�V}�<>�*6�7���ɂ�Pg�@e��cLVs�������7��P�\������g��"0}E�3Ց�||�+Kr�H�4x�ks�3�}ܻ�/
5ԘE�o�P�9����ՉIв�&Y-	���|��pz-���Gd«�2���u<C����$�N*�3�`����έDZ�?�!dF.i6H�̪y������6m�1O,OO��<A����ie�hV�T}En����.vj�عN!A�Y���o[k�R��L}<T��WT�����R�o��.���6�E!���	���zg*(׵2;�4�!�'�.Lm�A92j�����-���"��eq��1��x�o�0WXp �f{HV��-az/�H�Om�u��Ͻ	�����t�d�W���Vo��G�5ey���])0�hK��S@�g��� Z𙽫SI����ﳾ���Ȭ��^�
���ZF������X���� nt��Y&�f�T��:
FL^���.�jN�\�9;7�x+�q���q�����Y���s4����qqo�RL�I񠼱����XO��g��,�B_v�'��~����Ǜ�r�ړ�|�m�v)��+T}�v����`䷄���.� ����k���.ḻ��H�)��&yI�E�ǡ�F	m��Ui��f��78�$�?�γ�W�,�v��LX�)cx�q.�~����4G�T��K�u��3���N����I��Z�ĉu)bċ�!/������1c?a��.��_c��W�_�Y\]J8�{��V�h�l��(�n�����_�\]\���7>�GsG����Qs�!=��FZ7�I�2}�0RB�V7��峠ȕ���]�h��j٠5��L@*���jͱ�cᖱu���[bw+q?e8p3�un痪!�O]��N�g��/Qo^�Ѣ�q��Q�Ԁ�����QV�^M������o�������,vT%rq��8�#�a?l��~]Y�#���wߜf�o���I��v)|/Jд�i'��������[E��Aw�7l5)f��xoΠ�5U攔�5�b�gڸ4�[4��8ot�fR��2���L���+���G�w���E�`�R��p�����?�蒆G/�{.%����\�ŽJ �#���L�d���$�G���M����t��(�r�xj�5;?P*�
���d0��y�?���WH��r,x���ڂr)�nr7�{�&�#3���"#�rr3���$WT~�x�E�m���Dy �<�+B.?�d]t��.��C�N��R�a������mu�+�+C+)�+c\0&_����,�� 4��)�l�H�ǠQMby��Ip���铝���g�)�6�5���,�Q��Y�_7���v)��O**�F9���d���=fsy�Q8�Ld�-4���*"�� 2h^��bI����?@�(�H�@}:���!�K4��.�U�h�����
Z�ē��7�7�3j%~�Վ⻠+�����L�+���̫�n�[�=�oP�� ��F�~3�}��~l{��:}����_�C-��}�����h"��f�5d��M��i'`��X�k�ѣ���'�.B~�H�u*���`���G��$�K}Ϣ44��ʿw(�:M%��߷`�C�9��Y�y	ǈ�.�I�icȇ�0�+)���}��FPI��X�I�A�1�=q�q��jI��|�M��6;���ֆ��R�<lб\�����Wh<��&��@_�L5��l����ژ#�A�qc�0���MkZQDږ�Y!+NfVQk+
�FkelQ9k�}Vh)k��;e'E������Q0Q��<25�����������8��P�Yp�q!%5�O(М!z?����� ,�z�^���/��$���Ҡ%q;S���(:��Qn+����[|}��)y��H����'!��7ƾ�h�/�/l8�D���E
�@�΂Z{c�� ��
�}؅�����/y���ׯ9���'FZ>~��pz;Yg�����"��,Y�7W�Dw��#@;�sB*�Ks�%����ݫ����[����[�Ȑ�[�3Xb<���ɛj������{���S�6�/U9&{{{��S	�Q���(��/��17�+뱋I��o�k�4�����{9^Y§����Iq�`��F�+�u	խC]w�Um�,��5�R��!~%e�����HSź�W���]3V�����H��'_��9Hj-|2�>���J��� �
H^.�����sS��Ջ'�k+�����r�ħ��=_X{�d(D��Z|[��2�[u�����U% �+ԄO����R��\��/��a�|��������bV��T�"�~���"�ȩ�-��u~�诘u��h��*�b�R�/b"�n}sFa'�X&:z�2�ީ�2��i�իC�>HiK��_��c���_�LK��Rh�5z�z-�C��A���Ga���j��.�+Ѧ
&5�ٚ�DHt�W�?�x�ɘ} ��>����ILG�=���bhI�֮����;1?�2����,��3�,Bn�x*g���(s��8��Ei��PGhh8Y��Z@�r�B��b���2���gcǏ�oE���q�/>��e"��sl��CNO���_�vS�tcVԼ�U��ퟮB����@j*����3�&�v7T�:���X]���n��}A�$�2�1RY�<��F/�	��o�(.�J�;����41�����~���]�)����+�#��}8<���b�����-�Iw^��U	z������2H�[��� �IW��ېʩ�hk�D�G@Mu�<���[{��$����0`��~��Q����N�H�hW��I�+F���7|��KF��6�W]|�֖�u��q��S?>5��61�i� ���1��O��>Z�_�]�=�=����f��C� ��2Q ���Nz���$+�������:F�of��ɋӞ=��5�'��	��g�/Ƞ��~i@�/͗j��Wo������[*�^�-k|9�yR��"Zom(�ױ� ���#�ʄ�3N^�tx!���8^�{ن��	E�0���C��+�1;�Q��H��(k�Ў��ʻmz����S섅���%�IW�t��l	A�.�T������?�y��v���5ƭ��')e3sʖ�O6$�Vnn����� ��Z�  �/̜5���ޣu9VM���4�æF�:'��!Z��ױ]F[E��	����b��k>��hr~��%[??[�p%UggΦ����� )0R�k���|�6���ؙ����W���2�5�k����]p"����`E�m�|s�3Yw���IfA��� ���W�Y��s�/���*�V!�U���+_�>�	�u�뿍q&y0sY��f������O�����˼�4����V^[����7H��Jg�'���~�����v��Tar}�0�f�}���Tn���R�WE����+[� @ISS�[�O���I555A*#�؛.3a))u�@���s}@��,+5s�j���n��Z���E�5^S��f���F0·��`�RM�h�5K�;w�S�W���B���0�66^x�u wG@Hhr��}ࣧI��7b;s�?h�ٍFH\�}����E�q��|sBeeA�9��/���C<������צ.L���� m ӓ%�-�<�O��{��ehFW�Ā�R,[���l�%���a��;�z�)9����)m�|����"��M�����h��{��^�Z�񡡨���n&-%[a�L��0��1�;g�`Sy��m�_k5�e�o��o�]"��J~WgD�'��g?�v��>_��rв�S�K�s�����t*A��O�oyf�oG�C�<��얽�= ����ߟ~�ՌT���3�uȩhlζ���Aв�c>��G��UӰ���Y����ֳ��R�Z�?Hک��YPRQ=���Q#��
G��5��ϟ(@�i��*O����~-�IaZ�gi��&q��0��fR�����IQN2_�hP��_���%:��1K7�nn��F�
��E�333�::a6��//C Q�K�[�
[c f�f��u��8��J���y��/Wx�]�#��o�L��fv�k��E��H�YW�B�k�BQ�J�c2��}��J���q� 2�G|⛆y��"��^2m ��~i� X֓�P�R~��IaYh�fOv�Z �����6����ٌ�v�J_����)D�?��@׎�c޾�)NG����H��)�<RRR�N챲����ǳ��yy�hh�Mtu�&+��z�ǧ!x[�H$�DU�/R��U"|��!/���uе$�r6�*����} ��		��|�UO���R��SS=�	T�{{E��t}<~;?�s�����F�wñ��L�j�C��ă�g�l�9�y*�陪�ðk��U)��8�<rJ�Q}-�be�b$'")))���7�L*��L*��^o��
{��r���8�����m=������Y��=K�4��Ο;Z���8�/�d$�>7�����|���oY/OWĪ���������8�&((�^�����ϯ��M}�%Z�?P7lA��<Z][�_mCv,��n�z�[`!���+W�C(��nDgb"����(��?�o��L\���MNdH����1�j�9'0�ky�2mnd��[�J	��3z�a%c^l����㛴
u����4�S��׍����ɺ�U5"��������ULU���O��֢��
+3�U������-�t��s�B:::�jj�`ؔ7ʹ��Y���6�2pN�Y0j
��X����Z�� 7���+2��A��:�y�������}�������($�<�T�!��	�
���Xn��������f��e4/����W@��	@z�I��;����s�)D�(j�>��w����}��$�rK8fkw�+C�l�ݗ��ŁWRPp���Qŵ���3:���%W~11e+�P��P�����x��;Rot<�N'FJ���F���Hr��	�^k5M�>�Q���-�$,,,�99�3:��'�rZ&&&^9.��ɭj��l�����&#��S�S���%����� )���o�[�Й��i����� �<��*G����d���"V��7D1o�n"J���䇉�&�eAٹ5\�D��.'?�49���Hi0�W�~�M�����1�=8ؓJ�Uף���9�d%F?�aKfVVQ�3�Z�W��v3<� ?oT���Zhj>�c׏^\�9�]$�0�,�ϨD�����#->�E�:,7`���<����Q���_;��,[H���k�;�RD�t#D�O���u��͢�A�w��$���@�oeA$�I!�{{lES���aIU^+���·����������-nχ;x#�EP��7��6��v�-J'A��Aף@)��=�kY����f����/���s"g,��M��;�HٌP�ah��gd7��{�?�EބE �H�8���K(�EE�F�ήN6���W"���1��܍��Φ
���;X��'bƶ斁8j��4�m����"����ȥ�9��3��]gY�~��W����x}��@���*?�A**���X�q�2�hec��\p�J���
]h�`�?-9�k������#����X��JbU��ٲNI�"ڜ8g���K��P��x(&~����#�����9�~y��3�c�(��$�pTݒ��7�45(�<��=�e�{uW�@`"�Cn�ԜHb���%{ޗpO�v��޶�9Zn�<����� =n}s8����W�/~�]�qH@Fs���<`�R��|��A�@F��I��{эK̥��I+�r\`p���W>�/���oxzp��d�d�2/��!�~y?o�[T��>�Ռ�f=��k�0�YI׆���9�l��^��j�ٴn�|����1
]�֔"]�{{e%�}C�k%���D
E.? {!a{(��[�
*�]<7�`��=�:4,� ��n��Ϲ2}9t2����T�ٯ��V8�.�p��W�e�j	�O���vf*N�F��IMަ�=�[/����		h��VU���mۧ����QrR��Ze�^4�J�2䉟=ky$ ��o�Յ>�Z ��7�)��Ձu}��yf�pc��>u��m�533��q��3�e��Ī�2�\��ɯ�P*���s�g�����~ѫ�X2���n5kl��J���a�j$2v���;e���C�l�N��m�m3�ļc++��\+���D��y��=��#F;����3��/��8�n��H��|�ݾ�;���9t-�@t�x��t�����rr��l� ���kGR�/���Ɩ;��W��-���rn!�E�^>>�����S:���;=�9W�)�Ii�'�˱�+��;ͱ]t�;����mn;}��a�g�LN���е���sm����ޏS9�~�|N��=Kp��H�=xGD������2Y���V�}y���x_����n�;���J~(��c�k��=y3`m�)2bu ���g6�H��J���~�/�<?Ҫ����y�df5��R@X�/u��"���agT[�te�v�Wo��@i���ٛۓd�su.'�F�J��DU����Mc�����환�����`?����=<xGm�\3�c܂jӏ�aQ�4��ԗG���ь��o;�q����������u5FE2�����%�GOJ�q���;�-D �ijeE����	�������P�Zj��H��[�����S��U���-�<b&����G�hq��y�����CYA
����~��{��Ի�kX�Dn�r[�IY��߮�Ʈc��"F����Hy����� �(n�k|^�#�W�^#�?����Lp�	H�o�ⲅ̯���	�O��GҊ�<��w|l���^+S^uI��ɍ&�^�E��J>�QWW;s�@�ѣ����ϨmU屣l�];�XX�GG�H���P;���I�|�d�<��qJ]��#������TH���5>�mE���X�9k��2;x��gI�$��ό�B�3;
  h9��2Dr,� $V��n�ZP�9?(�WNq.7��m۟7�V 93Vy��<�-w3ԝk+*Z�k�fe���BwI.�g^'�����ԕ�yw�$��d�~���uVd�Ë�&��.�֢c�o6�˺�~IW��v'�:�k�Ek��o��Bܨ�JU��n�� ��^��?��%D�n�_w�;��b�۵��dټ�8a�]���%�0xf�����2��uJ"os�C([1��!1#���r��8a����rF�JKK{e7����wC�7��X]� f�==o�K�o���I���$ƣLW�y��fg}�)qJ�ɲ��:��)��k��2���^���{���>E%��@�_��>ib�䳘u����s|}w��cm�e!%''G-�-�_X�vqq��Aϓ���Ǻ���]���0�V�'�YJ�]L��M#�*v�7�&��� ڤ!��2#O���e�7WW_�}}F���Y��Xug[iџ��"i�\��$	��Z�^&f^��؇�و����)Hgބ<1�*y�G17��3�]��$]a��oɫjF'����JD-�r}[;�T�����
H��6?L/��8��y䏟�T���-��H1�I���.�JK�26������,�5�\x�QR_�|t���F��\��1ɱX��s�}��{{�Q�Y�<N�8�����d�ІɈ�� �M�tK�`�R^@l���U@~?�l_�~F)��BG$,�v�lL�bo�Թ��?̧��
�4*�S���|:��E�:���!��2-���jGdhB�_�}��"�|��%ڙ!_�=855��l'�+�GM�1�>�o�t[�gm55�K��G$�W��l8YI����cN�;Z��U��D����ʴpĭ�Y���Ko,/* ���#������!�,�R'�`ɡT���_�ҋ#�f@�����`t��F1������ZW��V���]a�ӽ���M4nnn[�7�M���g��)X�'�Ň(����A��VJu_�@�7k�D���ߗ/����䍡�i�����<��������!ggk������,,�J�#HުMG�}��X���������s�����`�p�/eR4U<����+$�2�@L�Ҭ��=�B9�[���Ȍ5l��m�Ǽ&LI�5*���M�{�U�����?K6�u��'��;��U��e:k�YӲ5�A��/^["�mHFL���g����ٺ&"�#����Rg�Л����ǫP���1�:&[���k���9��WE�'���ƭA��O�_�)Q�.C�f�|���  y�AK>S��!���3	�����c�%�2h�
�'z˜����YYY��D1�i��i:LLLнĮ�!�B�}^2�(v�`��#Yx�{��]�j�!'ddAR�\����w3����8���v3����>d�G�`�HS���4U��6p87uZ!��㛅��7�)���·��^
��4(�!g�S�U��f%7�����Po-e�����H���:o��0�Vpi�sp��ī�Յ̠M˿`cgo�_Q�k� 7����R�ʍ�߁���]\�8�d���Z��s�+�(�MS��<�7��sM�1�*��Aˌl�Bn����ai��<w+~�d��Y�)I/���"������![  ���U���U�F]��?����|�{|@���"���ɲ0,Sߴ^Q��Τp@Q��N��3)Wj3M<�a�R2Φ����w�.� �@CEa{�tY���l� �������\棋,X�!�D������G�R��b\�L��6�Y;ɲ���>�O�mvT�?��M�{�����*iL�~��<Fy�xD�Ƅf>�6�D��������P=�F��|�ڋ7O?H��8�h�6���4�04A����WpVTu��Z&`��ZF��N]-ت'XK�w���������_�Hƿ*����>)�ז��UW����x'�84���դ9����� ?%�G�5�X3��B�>���1k>�/�y�[��'@��*	��fZl���NK#c�MU�z�L�b�:�,)j�\��&W髋W)Ò�mYND�aX�y�Q��>�.�z&��8,Z@�ݦ����-]M;o�G�`�ӲM;Iǚ���S�U�C������1{�A�������z]���� *!]�1�nBc����fÕ&��bcA��m���j�h�n�'C�5#Ħ㋸�,��c�	*5٪|7�T����;�S΂)
�t�����n���}�V�}���"e9�@��3���JV󵘆{T+��\� ɂ	B�Ǘ�p��!v����&=��QhX��⇣�3=��d�]�xxԚq#��֘�]=M�8�(�d���������Y���eI��0�.Y�h�l;n"%��\�FE ?�>�"?4��!VÐAy�1�s������O��$��q�75���vϿ�Ko�D:,���x���V�X�zc��%x����í]��F� �]?�Z�O#�VS��Q���;T5�������:�}�S<Jk�u$��iT�'����'M�Q�t�b2��� n�����j��� �����W@5�~��� !)���t���J	H�t��ii]CFwL$&�F��Q#����?�sx���3���>�s���<�����i�-��b4T�<���b��IV�:�m�f���l��g�]�2�pߦ_K΃f۟̎|,�����s���j����M���!�&#�t*�De�{[����Q�
$IS��M��&��������a���.�:���i.JGA�Y{s��"ߘ��j�hJg�.�h��4*��� ~;2)k��v�;�Z���UU�+|��XPj�}�2}�s+2��߀]��"���B[	�k���mp�L2�o�/k�[b�D֒%:H'��?����D�c_Ϟ��k0?�����D��q������h/fr֔�ڠ��ikb67mdrjhh�6iW !����}��S�����.4T
�o���y�{�k�#���?�F�3zX�n�N~��dV�Ջ���mE��<�L�l{����]�:�4�K4��RIl�d�A8�b��q�����z��(*��%憘��RJK!r�G�tc�'"��bˇ"�n���/I��!�'�@�����J��S�����*mW|XU:1ow�Z'E��)��14�׼10ks�P����6/��Q�$�)~���'�;|�_|%���9(���R�OG��P*�,o�4��ώİ��21�m\�K�����%:>ש�RI����=?��� TdI��y�6��0*&�����Ͼ��`^�_7(~�3����������+��"��A{z�mm�&ڒG��<���x3�S2���
�U~��6�w��b�ˤ{V��P�&�P�}�T�퀕�`��R�V�R�O���5z
!հ�Ci{Z���:)�Zi�������r�G�G�/���>�c�a��[I��<��Q�[����d�A�rYrv/..�a�4������T�0��?.�
�V���w8�6|�~��P�t�e$�Xi����6J0��h���[��3���"�7�,Z������J-���[��o !�p� +]��5��u��=����G�R�v��V9F_�D�ޜ@6�;�����:���C��/څn�u8(k2��܍s2s��<󶶶V�t��m�u/B��3ֻ�����ᇿK� ��:7ۏ���;MtX :i��r{�w��x����@n���R`l��2z�;���DϷؠ'��J���#1t!s�=M�o��C��*to������By]#m���|�`J�la�䨮�%of��C����.yV,���|U�
�Ѝ��Y�gs�P�����Ҫ����{Fx1���P�v��=%5�r�f���������U&�m�._�Fp4���Yc7	������[�.8��r�|3���c�����+|��|��9v����~1��fw��\,mq�$����b��SО�{��[�W�w�{V�7�U�{57��߀�����o#yw��nKП�:���I�����X���v��$��L��Z ո̪�-ET%[��+���F�y�>3�n�4�X@���<�b���O��x¼�<jyyx^����~(yvf�C��m�0�)�Q>������ן`��p�����?��uВO.}�#涴vE��!�zm$��h�u�Ե�7U)���Ue�ˊ�$���aC`t���Nꩃ������K��m{�rS��[�|}/��#�UHD՘}SDbVqp��������iJV1��ʎ�A0����I��NPC%�27��ê0����X����쬢� �������F��X٧��3!���������;�\��1jta������!�Ū�$ybi+�M߳��v�`�=�jB�X�l����{RjN�k�C���c�?�^AGxtϐG}]��,�Gd?[rʘ\�E6;���@[MDU�H���~�w�;�7S�V��YR������#(�q��������3��R����M�Ix��_�B�t��$��fsJ�!Y�3E�T�I@��$@����\�v�#�Bxd�A�+F"Jj�B;���ĝ��[��{�����%�������w��TI��mBY�릲��_k����5��ƽ���Е/�\�;u�!�z!Typ� @"H�w�I_t1�-ϑa��卲��4=�36��`F6:�cqg���:=�<m����1��`��{�(�[��:�O�Z��B��y*?���"I����Z�P��|pPõ�,�xH�O�B�^ʩY�]����<�s�V��+nhH9==]Vrnniygdv��� n�x&6J����.͛�/�\��*�n�IGmz�(�����P}�~����=��'e��$t*E٢B�?�0�~C
�[>���gz|峲��'%%��Z��[�GE�B�4��Yg���Z�+	���Ǌ�%"�|��k���n�Ig5�tV
�F�^�i�W>�d
AKd`CPK����hHV	}_)w�j�<��209^����ݤ-�{j�Ϟ�O��.��Fgb[7[&�B[�'����ɀ���
x�l�r����{�e͹_�4���ڂ��Z�z�~��%�#��2S�aϢ�һ���~r��0��=ox.`�����ۭ�����Z���Rz���5Y��?n�"Y�}�9؅��l�@%a�����=x��y3n�rC����Gۻ�ĩ���~�ٍۚ+"�ێ�=�����j����6Ţ�顭x�!R����1��U�WW����&�8Tb��>��;0�H3ٽ���#�{鎉 -�/ׅ��Dk���C��]�~�<L�(��,�0\z.�Va�W?@�rdGo\YU��2��Eijv�_���#�I��S�i��V�9z�A�/%<�E5p�S��Og��K1��;�3�8�0�)6*gr&~ddGy�H���_B0ۃ�Vq`z�����Х�6=9}܊q#095R�\���W�f�i��`n��T`�@׊�z�~���p�q�����}�vp�k��L�Y|&\��K�iŭ��z��1����bּ�zqk�(2)T��ɬ���u���9_WP�(".M�3�Yh�kk�͇�i8����x�Z�9����@�'�.���t���������Ց2�>����,H���`7O�A�5]�d����܃��^KCѩ�g9(�pҐ`�xV�_+����0��Hȹ\�V�ģ'@ �; �=�(Fj�	��*��������7�
�V(N�x:�	WI�Vv�k01�G�,���+�?�>��:H����$F��|q�˗F=�����"�Cf�y#������q��4���ğO$���,���v�\(T�
�s� � ++�A���h�a�4�ǎB�÷�X��zS�Ґ��5V$�E.��g}-dnn1@Qe#��/�|��I���� �y��h��O�J��.������?�vu@u�^��~t���3��܏�C��ۧ������D�_8�U�j ۝g�F����(�q�{v�?�$�=��QX�`���0��LZj�"
��X�p��o}J]Z�M$"�'�VdzL#�E[qs3䏂�f���SW�C�P����4�y�gW�x���V�Յ�l1 ��y��{�^strrr�1����Xn��5��4wEG��4qzI��n�x�iht>Q���5J�Q�0/ϴ��gm<`�7/Dhj<o>�J5�$���<Pi^�"|���{��(a�7������iJ�$������F���F���Qf1W��I8��O���skF<o���x��r'[Ë��le��Dm@*L9�pV�U[^e�~��+��r�8��4F�܆���Q(q�L�؍_������|+�'��#���ˊ�0d���]���P��|�&.C1�EN53Z �>ꥤ�oB�Ĳj.�m������7'��ŉ�����Ϻ��ז0���c��9���uEYي�7	&~�H��-�2��xj~ߍ48��Y<N�QRR�:���D���y���z-[�nf��"�}����9�WҬ�����?~�7tS��t��>��<�4Y�U3e�u*�� 4���<��y��C����OZ���c���2e��Es����a����A?��*̓n���T©~�s3f��1C�xEV4(ͥ0^^�l�r��W�瓐�O~��7p�3c�v��!�����^Qq���"�97�P�l�q?�<O%�ե��k��	!��M~�ߖ/�9��cZ��Si��S�V2�v����{� �����a=��EY�<r��b o�'ql��(঩9�`������y��p��`�tdA��0L������ó��)�zg�ǉ���m���eo�#�
Fm���pgfgm��`�_":?=MO'�7�=J�Emmm�54P���3�4ү����y��$q��(�Ѽ���.6���?��ğ���h�g�:�����9���\��x�{��t�7�d�0��nJ�9����96Qa���3FF���ڡ��!�r�����)\��{b0��ͨ�����u�0s��`Hb��e1x�t0�#�hrΥǘejA^S�9�>yppp�(�:<�������!wâ��d�7�m:w�^ah�6d�������`b����2�}��`�5U�/����sy!�s�C-$02ך�`�y�M#��T�BB��o�:�����_O�f��vq�v*�������t��ط�n>E�y�gW�k��)OZ�������������-E�{}~R�zd	���?��vPѱ���T9����*T�?1�����n��9��sݘ�� #�t�c��涴d 0mm%l�-�L|�DII���"y~�I�"�r=VvRp�Dѷ�熫aG0˚L)�d��W�~��O�_J��Ofe��z�v/�-�ɫt~�{��|M�F%ZįLu+D���vS�嫱@.4�ѝ�:X�"JHaH�iz�U�����'�'l�0�U�'D�)*eEh,��(�_����~�
ޣ���ⓤ�B��ʕ�M�~A��_��&��ϱ�{u4�T�=*��m��P�U�`{cg�qrr�qq4a��g���N����w�}.y���%��H�yU&����6��p9^R��
%���F���j3�����������-�X�(Cl�ں�Bsqy���E ,���j���U��]��������r��	f���K���D-ܶ�H�ı��T��"��:�2{ug��s��v:��9�f89]�΁a�ǆ����N0$��
4J���C
��R���^�J��v�/'.o͜���9DQ�;���%���ݡ$�$�d/_E�;3$�t�	���� ��mo�S���>į\
��x�gT������Y����Q���8�'%���-	��Q]<2������,��q$�*�6Soll�a�1��=�lvꎦ�`٘�8��_�@�z�t�L����6��\4e�:�S�W�Z���eX[�����v���ZBCth�m�dYE/����Zse�X?��n�@� �����!�������S@�
ߟ����N�H;�7%���0③�.h
�N�n>>=�m��oYW��)���c����uLL���S�x%Y�4΁��δT4O�fh@a��96i��Fb��г'�Wd$Roϵɺ�#o^d����<��-Q`x���q?��f#(9�&_���Gt��v�qfF� ������0���~aٕT�?u�87cb���|�7����l����n�������a���/+"����dy(3��޷`����.�z�p>�q�P,ְsi���K�P��xL�=������B&��c�����d�۸�!�ްrQ%q�SI�A/@�P�)5���C�����=�^3ש`[9��3UxGw4v&��I�	�)���~�����L� 7L0[���T����7�>ap��F��0D~[ۭr�o��*S��ⵙ��,]s���~nM�L��蝋c4�8���8�̗��wr�9�s��^��)b��蟶�$('���Ty� u�Z$��r�p���$���r��ٚ�gOG�N�#���j,�zp�_Q|�Sb�ͻC�K;�c/�����>N������'$0r`���D���=lB�SPQ�vk�7]���ޖ�Y�����.�7��U�@�g%�.�!���WR��i,�aw�,�`-��y�������HJ�I*�t�*1�����4|d���W���A؜djn�0��u�h����?_����]���CY��޲PQ�uQ|y���L�%2��`��b�6��ſ*���1�gD%�e*)+-*,�~�#���'7Ϥ���;`��h%�E���$'>p�P��P�j ��d8>/���c`�x�M�������(�x]�A�s�`h�9¹{gFO���ԠW�2���e%����g
q4+�����/�>=����Fq0��\���g[\�����+8	�h�U7ԍ�D��*7+J2��Ί�$�=�IT���Ϋ4�Q�W>�<$�Z>K���$��ݿ�<D!)|��iD�٭(������BÞ�ة�V�"�y���̓5���wƳ�qn��{�nP�J�����De�2Z�N@�~���z����Ǳ�PM�ZV�6����y���r�~Ԗ�`T�|W�Ȁ�.*�,V���1x;z��{����2�a��ӛ���+�{���7��?3�,V詓����k�\���X���ee��򆦦^1$��2��wk&�i։S�}%ۦ�_S�Ա%m�>��o&������f�,.���@� �J)����^3��ܯ�"�ϝ'3��-��ԼX��㈒14���s�����m���\n���P�bb��vvv��V��5P-�c���i���7v��R�7�+�O�҃M[	
���K��K9¡;��L��2��)�-7F�7��?�Wʰ�H+�^5�VsE� �ެ�h��J��{�*J�tt��x����G)���=~aGg��}Ĳ�սA+..��ч���vIz2-�+�t��?���P���%��YO�]�n�dJ����\���%cc>�cNܝD��+���5�z�td����� �y�B7�/�km�w�j�wbx��DJ���Co�Ӟ�:k�����V%�/6B��J�*�\b��Bk׾��������#,��;-���k�,u��>&�y5�J�899n�����6�h�t��=��U��|�R��;&x��N�X����s���T�?IyH*�!���MV�u���w����;��S��HvBD���266�m�ܡN����M����e���Ӿwm4q�T}�I�.�Wמ�<[ƥ�X��%aw{�Z��H̠�ϻ硂��s�<Z��a��_l���?�����m��b�K0���������%7�(^���{��f�Wkd&�`��������Jl�$�,��I*;AITH[ר�w�i�{�A���kڐ�p����ּ�s�GwѮ�����՜�U����j�[#��4��3݌���	O�2`���|����:uWU��-�?�.�K����v��=U��8Y�v���
��u�T�$��6��9�?��̛e�a(ޤG]hh[w
x����H�\� ;�Y�3z�s�ì���C�;R�K�<Y_�~��]�\��)�H�$�l���p�T��g�KEf�M�I#~��U����-����

TTTKW($b��wk�b�>���B?������o7�����\[�!o�������ieD8X߭9��f�h�&7����_��)��ٞZ�8 [����g�Kbt��K�t�+IG���B���J��\hø�2j�������T%5�G�BJ�֡��W�9D���zRS l�<�EIM@`��v
z%%����-����­�g�gm���X�|ozzW�#R.f�:��mY�h1+� �Fؑ��lv<lz8��(�-������~�t	{o(���QXA��:V��,/�Ï�̱�t
5�/=&-���Q��g� ��B���Q�x���*�Cz�i5#�Ƭ�۫�DB��LbUY�-
	���T�S&l߳~9��=��B��2�bL�us��_��g�:6PHHȶ\�l���ϥi~���ԫ�����닙ɍ�}�������������7n뢷��$]��}_�� �҈�"�/�q�_��rN�Xi�J��s�l�n��G-�]&�Lb{�������0�x�＿�
�W}֊w�7o���tZ��c��!�q(�]-wb>�h�]w��]�ӓyO�� Vo�+ӝ�%86��Y�g?�%���x(����8p+���Wr��g�:&�������@4	��Y�IJgA�?U�����6골�9��ӣz�����s��.W7�7�ž?��ī��Y5��XsoBVGU�=vZ�/7��e�?�/������7�P��Q�E�I���D��Q����M�?Df!4o�_��_f���5>z�O0���PP�����L`�p]�ܯdZq�O��G�n��n6��0����/�#���s�4��cOϨ������g�}3�71� ����n�5Bڪ��B��=��%]�8���3\#'��i���V0$f��ĸ�����?��/�QV���_�t���/=9\��
��3�.�P(���s�U���z(=�o�����v���gf����{��'ϗU鋸t��ϵ�|�,q�i�s�|b�	�5��o��=�{�� H�7��q6͚�z�7���S��T��:;6G���[Uq�֜Ώ)���C5��m����ԣ�rw�a�9O�hˊ�װy�����>&/
���Ϟݭ����U-|��4�R߄�ҏU���s�m��/q�
��qDf�͵�z%/Lq��T��fY{������L�d�,&�
v�2U5S���i+Sװ��9s�/c��F����d��ً��$���I���}��n�ߘ��'8�����L�{P^q���6v&oh7P����z-�g�_v4x�I�>|P�I�p]���� ���C�3�̗�so�g�Ƨwq�F��Ci���M�7D�¥R>5��=C�֪�P�>��:��/Q�:$x���1��v�����^��wᏚ��������T4��:���**�7M�L1ˤf�7��Y����^�L�n�Bk�q%Ά�r����r�����s>��T���Z	�L�,V3Q�iS����8�ۅ�'ꭡڞ�!�Z��Zn����Mbr��_��f{ph2�X`w�B�7Z����{���?�}y��N��dQ���m��A�;������G����_��2��̈�����%!��R�����I�����syH��OD,6Mk6%m���,s�r�$�Vi�p��c�)����g X[ǽ�^Dճ��>��@��OQ���i~|��m�(&$�*4W��%P�{��X�-��P�C��u�Dm�� �E�4�R>�^�i�a�r��sa���w�7h���ʂ����L���Rfq$���lb�S�"H��se0�r�j� ��؈���ز��)_�ؙ,�s�_��q�6�h���};U4��T/c����z��9SG��Er`�NC̓�"�YwLĊ?�i�<��N��Ϧz=�KU��W�=p�-0+�h����~��xtjWP���C���KO;�tJ⧶����ό}�L���r�(u���BO��r��~A�MZ��Gg�&����?d�~�&XP������3C*9�pX,������;]��u�K����)�:�=����>�]��Q0��1E���R�̯Y��Ƞ��j~�Y��"��P�����P�ҽ��G���BfY���(,�X�q[/�>�%{m�'O�%=D7��Br����3b}��Nz��'O�/�w�h׮��-r7��!��de{:���jܲH��Kz�*~��?ٷ��[T�G��Q;�pQ@}t���3�+a=�)����x�
�r_Ս�͝�䙙��;?���|Sվ�g.��_�a��X���9d<���@��pIC`~�k����#K��dL
Pf�����&�d�p��%��٧p;FA������lm�j�2R��`�,�ʬ������^M��(�����韬56w��}�����&ѐ���em��nD�N��z�'��w��I��O冉H^���]c�0k��>>�*�b!��Zs�F%꟝�������M��XO����ı��sm�[����@Qyl^@���hn��������6��(�b7�\��G�-�_m|�6��HÀR���f�w+���Kc��OT)v��0l������tZqy�z���4$~s�LL�=;�߾��{?"@����P���}��g�g��&1�%(��.D�IU;�w2RU��t`Ԫ5E��|j�k�"!Y�Tv0�شΣ���Ӥ�������e�)�^��7���z�v��i�����~���4z�\�	�s��FG��*B<R��������+���j�o��!{�:�}Խ�|;����O���KgO���|	�RU#e�C,�5��=�Iu5[������Y��-�������ʉ9�_�azh5���2}]s��(����~I��,�<k>-��x)�B���xE�)�&s��kѢFI���'�F��<�t)�ᤕg=�*zr�W3y+���Q
����t�Mq��X��h�	��I��Ic�ʚ��@�V���R��Ќ��R�f‑ѧ��j]N#]��d%���� !s�@���I���1{��u.��f�Ѫh��q�*���~��5�]O�t�'4����ղ�Scï;i��ℕMx�>{�J, ���Bc0���Ȧ�m��3��[m����ch��ŕŉ�RK&I0u�-���\#e~KѹӴ����C��)�muU[�[&	���gL�Ȉ��QQ b��g����)�}:���0����\'J?����'i����ȕ>Ǯ����(����]��]`H��L?.��W���ʱ���c�Ee-)����a����T����4}~?�������f�����ȉ̊��1���F1�v��pG,NV,��ݐ/����kO�O�S�J���h�cZ���� �(���Ɲ�U6��#��)��^�r���yG�������$oh�g��[��5�M�4��#���3Ku�8��o���Ωze��K��s�t�߰�����͛���)�rk���ffY(kL7Ve�577�ʅ����[��붦ff�xzơd^D����Ǩ/���U���Ճk�Ԑ������/Ε��������r�t���u��6~Cx���	�+*�	��ZTUU�$�j=��r���l�7R/����&��+R�x����i��,��2���)55�ɜ��{���cF�V�@�e�=�t�rF?�iJ����0�ϒy	���1)���8�ڿ���#�Yerh�鄎�D�u����0�- ,<:7�\]]O�{2�*/���E�:�IJJbfï%�yo<�Qt������7��=�:G�ӆ�6��,ҕ�oHD��QF\Mi���<%%MAEE�3�J2��c�)1�-T�s�K�Ywʛ��M�2!!��m��ݐ�x"x�����)�_U}�Bx1ʄFe�H��\^���Z����zz
W���u�!7�)WMo�ҋ�,�, ;�	�Z��W�"���>��^g��7��Z��=[�M��K3_Nr�����@ee���᪁��q+Cc:�f���*@!�{f+9�jL����K����/��Az��+��*���x���)�}�ńŮ��0,.�[�3m��r~iidO��m�`�(M)|�8v���U�q�ˤ��S��>R������hO�Y�
���,��a��4��Q��ꥤ�F���!��@���޾(�:���W��J�a��(�H�.8b�M�_`f��ir����r��&G����MEA!)���zw��]gpK��Ȓs���%�~�h�ȯ Z�D��a��������򨵃Caa��0bqk@]]*ZZ���SW�������ஒ*T�u�2u�37E�����	M�M���+]����1�
^��$���羅iڣ�j>��96�?�E�����n��Q2ff�uuu�����v�� �ۉ�M��C�r��΢��cmE����@�7���w~��wp*��O�"�,����f.���>�]���y��ӧ�sJ�8w1��685������ó@�]uF߲�� 䘹�1��� ���U��3zxXʹ�����k���*0�=:Z\\,p�T��,�������������z}��|U:��z.H]^���U:�ևp��#Q��멅��J5b��G~nB��{�7�z�IR��I	'_������W�'�@����\�B_�O��n�7&&��f��x$�V��(~bI���$�P��<��t� �rW������K��yX���p�p��Yߡ����;n��j�}�L���s�(Њ�!�}���֖�8v��pma������%���~���>L��hY�A�����q��+m�У3H��YjE�O::�@��2�QE�C`&=%���p~�t��S.�����s移��T�K�n��ߞ�:��n<�4����{�(�޸���X���� uu��L�����^���tD����1���q��'r���S<v�Vx�+r�yOa4Fn�x�K٤Lκ٩N�d����IҢ���.��Gy}}���\و�ţs���
qt���7�H`êAE�C�%�(/h[l���u�ޞ��O -'G���T����`��Too"k�قo����N�dwY-O���:�P��]y}j��s�|��s�� ���SwCV�A�i�xd��U��7�@"�MLO���ٹp�ҋV|膫����z��E��ބX����wNͅ���D�W0�c���W���F���3d�v�BB�	�D\W�1����q� �;�V�w�s�`ߛ����p��h��~�n೟��~qyM�O�dx��'�����Z�j��7�e��n�v�^�������Q��#E틒�l�7�"����2�;��G?D;R;4M~��wј�� ��c�g��4��
U$(PPP@-��C��o|���{O*�0�J�S����JT�4���T6�G�!�%�Y:1h<z�.A�(����`�,>A��B�H(����˟?��|9����Ԯ�����+�b��P��B�Ӂ}�iv��1�����.���VO06�����ҏQ���K��OT1���mVE1Ifɑ[�ߪ1����/�R�ģ���_���FY��~� �X#| ����˚�!S����E�]H7̹�$�h0���0��DKuD������XY"������of����б��k�
ڸ�~���O<�%0�]oLx��u�8u��BS	I�A��"��۽z�T�]��~�s��@>�Y[�xRfL1�4^}^����˔`M5@�>5�y���\Y?����@�͚���2�^2������qחg����́���~�u��w%��*�."��ա���`�UIY&���q�W�ay�W�{%�tӞ��!���1�������~�!����R|��s~���9 �ܓ�r�h�\a�W��Ľ��A����&J�� ��%d����W��(�CE{X��"�l'���F�	kg��\{��Ff�ݦ��54����<~���� y{�]^^��fۼh�1@`BY84�y;X�)n'�{�C�J'��wO���ll<�nYx�G0�P�]P^�vf��2���l��-Fy��T�}%#''���Y��ۓ�2�=�el贫�(��9����3�4���Zb����]����ٓU1�$d*�l0�&�w��r�m-C����<ʣ̿�:���+v��
��VU�T+�2%�����,)���s@[�e�n�2K��*��nC7�rZ���W^����cۙk&?�&�|3Ue�����?��m�
Χ�m�[�K���˱�+���U�S�ʊC
ڶd�cߏ
`��D�g抎����D�8��f�'�ǹ���nq�if;y@�Z����r����|G^%|�>��T�r�f�}�P[r���ކ�Ç�63 |�}V��.a��4��ӝ���kd��i_�������i��!����U������� �%������=��7�oq�Z��� �!��z�7(������GZ��V������S�vmU�0��S*�=�lyD3�Y���}��z�p�>lp��~fI���;�)+�~:I���zϺ��ޟ���P�����X���"�u��]�d�PE��_��n��)+p�F�특,�{�4��[�����ca�S��u�����&���7r��>�F����ј?!]�~ǳ��X�v�O�nb4����ڛ̖�,^�Abg{��|i�}2�Ya���t�o��|�+��V4/.꽄o�G���|��#�ۈY��f�����8�"ϼz������r��,��dx���eASS*<���^嶞C�����4�M���ߜI�wF� �'��@P)8oC3���}%)\�5~_���J<?�B��c�q>Q��Yt�~H>� %�1Du	W�J��+Hɠ�I�$I��(�nՉD�U���&�r�J}s'�������B�Ӂa��Lm[�N���؟JI���$�I��
,������/{����"�-;� g�u���4]�����m���� *T��.�W�J����[�f�n��J�W���a���7�A�g������b��x�i�CqH��U�Dc��7�Nz�)˭��m���;$�&L���ds�bb�V���I���SYY���3Q�x��Z|OlX �Č�9`��� �͎)���i�'m�cT@l{y�!9[�ۛ��ť�@�8	���I��4������i;��Ū��f�5r�3r$;��g�R�8ۿ�䤥�w(������E��L� �(@���ox��w��r~����q�#IO�n��~�����>�ڬ�6A!E��V�M�{�#�`aX��F�gh�T�����ߕ��G���=�>�I��.���]\�Ɠ�����M[k�W��*����_�-5�z.`5��Ioư���L�VO��Qe���i08�JO���U�s��ɳ4�knӦ}H�N�g�	��/��B�W��S�_Nބz�I�(|��TD˃3�J|i�3OI�u_����	����@㉡��i�VΆ)��b,,<e3�?��KȁQ�����ett�kh\H���:Q����Ρ�Ł�>ǔ���.�s��.m[tJE�S1+4�I��s8����"����%�v�����ҩ��rl^Q�w��O���'x�F&�+H�Fl�UO�Î�4��Q������V[�G�m�_EC��"��M@��E!��GR��;���d��`�'9g�������e"�L��V�'��~D� &��A vyyykG[�>�*Ά����domCb3j=$Ά������Cp�s
۔�]֊y�v�|:MN��WA�Pk�?��*V������v:�7��t�q$%%}�א�:��rqto����L�51Ya]Ϙrl�X�2��;с�[1��"�&A�6VB��6,ii�6�� �o��y���t���Y����'ʅ18D}�/e�c�Q��0��t�e.�1�
+43xp�NOib5TqG� ��Ѳ�$��S����&	Z�^2�h��ij�s���ܔ���@:b|#�H�pO��Y��g������w��h�7ҽ*b.6H
%�+h��y&�j�ۮ~�#��|����w_2-�(�����>������HƳ�=����u������Q��GW�@��}��<��;�8�	ｵS��g�1����4�ճW>������:Ǳ�~"Lp�G{�bːH}YF.�+�i�O,K�x"�~l|��;Ӱ�7���ۻ�S��ָel��h��կ��h�����Pj	�k����T�T�&8F?Q+��:�ެ'��;�(����џw����B�$%���_��|��['�����ݔL��guSw�IqkR���<WK���{!��E���G=
F��&�E||������v�o"Us6�P�)�,,�3�2	
��~��/��t#��r��'�P��l^��h7���x��;�ُ���F"N�}`��Ã��S�W����|��F����s��9)Dtgw�����D5�cA��Q�N���~ő�����e�*�3|���4�?r����y�� 7���=��!E�o���ĸA��w��Ԁ��1:���X5	�L*�ܭ�K�߁
�t���/+`��mH9���S6	R���D�l��݇���	��%>����-*�<�e�^��}�?�����<���o���+HY�|�NxA����mH|/�����!f
z�2�����s����f��F�p�,WMc�Xf���`3�k�b=��x��M�b�n�=��!ah�+*�Qf���iV(neNԶ=�Ns��1���#9-89�_W��ځ_Ӣ8�+����s��l�~��6j`a�B��s��۾:o�J��]�l42��r%����H�%���S�'�?�LR��\d�w�����ZO��/c.�)����6�Oݔ9�)��$�5�p�Ϟ�^�ґ�=.��՛�C�$���o�t�ު��|꾡z�� K���Kؐ|�w��Ac�����,�F��|p�8M���=s�����{���!ÿc��A�W����~���T�ˍ��_-P�#�9�<ͼw���b����r�ܟ�;��8g�Dhlr0ാNr=
8�|k;~���z���U�C�Gy��}H`g�n���k#�;l���(�f��`Ȋ���5���^BlGc痗ǩ�^6KZU��e��'�N�������ױ�-ܲ�e�X�����oq*S����c�<x��Ic�&+�/Q텏��
���x{�p���T'$�hQBDｅ(х�{�wD�5��0�E�������F�#9�����zF���W{�^�Z����C�Iq_ݭ�~��|ms7VB~�H�{��U2$�  T�������UU4��w#8���8�H�5rt�S)��>����VI�Mz�Ą�����A���񂓀�13Y����q��o��[�d�����A�G>��o�x�� ��v� �9]��*����v].��j$�����kt�>-������f?��Mf!A,��N Z}JӃ�"�Ӷ餆W�y7EH�c�{cWPĲ-��I�"��@˟��HI�4��b���ǐ�9�T���QQ��H�E�
��VO�־����^B����gן2'��`�{Z�e����ۨ����{瀧�ߣB�-ﭕ������F�����a��B��.���E�_h�Ya(�j�:q���ն.dB���_��!NGz��}��O��+�h�/��o�����˵<sj��v�� ���F�Ǌa1�b�]����j�*�� �gZ���s���*{1�3�� ci�rt���;i����l2K�9���0��9f�����ge���~R,k���GR�/��ӡL%z`D�C���v�|v$@���Ӵ��2�Iw�26����#�(f�����&3b~���ػ��H���d��x�JM<�o��eo
��d���-C���>�S��_[���K�%J��+<�,(��4e�Nu~ -+�����1U�~���P������X�js�Y����o���B�8Z�;�Ԫʯ�|��63ie��5d�3���h;\�HII7�����F�̸�ȇA�+cn*:b�g�0��7��vlW��h��$g^��m������R���~�Reҳ�e��x�{�Z�1��,��)�9Xd��.c��	�����D[��s�'��oo_�����X�5�����\x��Ǽ���a��>��=	�+��Ba33���P!���E�)��T�tG�Ѱw��h�L�,��QI��7_csn���A�ŵ�p/.z��Js���r���"L������>�O�������0�DqJۉ+�5�};�2j�����@�X{D����~N���y΍�"e`0�����؜��iIZ�I8G@h�j`�{�NlxV����9y�m��­Hq�6��u�p����f��������*B�x`�o�������gn��6V��f�Z�LS��&��2��8�Y;�~Ǆ�g���V�����)��_�jԇwlN
V�87�����š~�_Á�}���iJ�ʶ�~���7��"M���� ���7��:-8�(�n��]Hri�OV���B�⮫MrNr�'�=9E2d��ξ A�Zf�pnZ��4[Ã�ϫ�R�M������w�s�d�?{��'.�|DU���&�(om��rf��[t�K�QR��K���X:a���������������>B��%5�	��&=|��j�0��a�<���J�W�j��a|v��
Q
:NNp.��{'q���lx�()�*�I���
<���К���C�Q�8|�'�yG�[�t�e����H�ʠ��hs��4��qv�m�%�M���FtA���)�o��]
�/w�DZb�uW�10�F�KIA1���O����iDj��㸹yث�uF�S�����3k32oSG�p�i��{I��ik��IL��j"�0�@�o#��L��ca����Η�|%_�T5>Ma"�a�yO+�����5���2��=N`/>VRQaO�=��P�j	t��(Z���dl����oDXr�Zzv�Ð���޵q�wg�W-x�v��`�=>.'rr��^+��߿���R�Kh#d�Ϋu �#�5�;�b6!�ڀ�r�6��]�tq��4^�_(�YحL�W���k�Q�/�8
6������t��R��1#��%��ڝd���&�;�ZO�#--�J�����ҍ��Ri����;e���B�Zo������Y]}�2�����:=�E�X�;�'E5���d7N�m�m�fW��tx�p�ï$K�)���Ͳ�3���a~��PGwKn{xE_O�C� ��1�W��Y6��_�̂Z_��b8�c�N����-H�ֹ�+y��:���I\��@���P��\D��g�qtu��9hEl�4��,p��<I�}�xן(GNA���M������fl�&�İ$##cmw~l⑍^t�Rh��trk��zp������� q+�LxjT=S��/Z�\կ�%޳�g1��E�G����!#�bq*��J```?�ʨYi���J̛��X ��x�}X_O�q#�_���K��k�[�
?������	tG��T!�����7��Rn0���z�7U�ĝ�Y�j�G4���<�����˻��ߒьݠcq�Bɷp~��	X���:����f�z��~r�@f�ޭ'@O�Q��,��Ћ�:��z�9%ǟ���jW�);�i���ٙf2�+�Ia��$ݛ�-���P���rՇP�?���ePUUU���������7&2'��%|��br����z�l�@�4=����17��ҭ�cj�qsEo�Q�
Z�Hĺ;ʤ��#�6#��3��,��
&�!.��B(�a)d�`����,t���c`�'��lΦ�dA����8��#�E{������woD�o2#���_��y3Ȇ��,����k�o�&#]��0�d��%�E�֮�	bu��|�tا�s��cUg v���j��:�=�[�ǳ�iA��z"-_5�۠�A��UceӺ�I�x��-�@ZZ&;LK��Qj�KU�Nem�F�����1�bY�Aqx8&�!�_�l�|�Ib\�'��x��8VAu�6��}A�x�O�4���mj7A������`lb�%�C��o��������K|�3b'qH��}���xSӲ`��SS��r�1mV���I���g���@������A��#�"̝B�D��;��-����]thhh�5��.✩)]�S�>j�^?'�����Nހ�ⷶ�� +�]mc�����td�t
�n�Q�?	��])���Zu�W��Ӽ��f���Q�c�q�	Ŷ����Ȝ�}s�緜�%����ˏ��r%'Y�bؠW\�TN�_z��$�
Z�zU:��M�N��Z�J^_*6���`�OV;h 
\�$��S6X-MZ����!fڔ��6�ٍ�\��l4��8�ks	�(W[�)�y�(��/�*�>6�j�֬ޛ��hG� �W3m������X��n��m�AR*�����wR���}A	�I:�
���J��x=2f�B�H����oї���c��wF��I;q}�?o��a��2�8�R��3�:��̡3���1�g�G�} �Z��P�;Z��d��Z�����kkg�P���tsİ�-7'g}�H���@DOv�=�/�G�i�{x�M��P熩���r��JXʀ�ȉ	-d�����}��Nx�@���|�B��a���j}�q�s�^IzxCzwH�:qn��}Wg��m������q��u�q���o�j�~E�"�N��|�;T��+��e�����q6��db\L|ڭv�X6{��77���Qu���*��`��;J��\����;U��Bn��z$�@?~�TIf��9{{�z!�[ GJp�U�o#����V���������^������:��_X}U�>bķd�]Ql@s��9��$�y��m�@�� M�mEH�V�ϖ��?T�ͱdA�<�"s��u����9/�<##���p�L����o��D��{������cY���x�}����h����C�Ȣa��@��ɩ�qF�1U�:굼�Qg��CK�+��+���xX�`�x���efϨ'���ѻJ�ЂZ�0Z��?#F�Z��X0�?$$[G�	B��{毹�.'��7a�=����D,���]��5�\��[<Y�1h�{6
x\��K�����n�Կ��T�H�����u��d(�)�W�$u�}��/��_�C�5W�=�)bk�`��o����ʰ�՛���I�����5��QXI%���[͇6���C�I�x�,+cO:7@�<�.�S]�x�vOE��@qڸ���3��.:�����[�|³���UW`�X��S͊k�s���nM��"�7f���i���<l'��tY�DFv��DyV2�O�UN�΃��sfp���i�WE��)�I�[lML�z���~\L>�}�|�X����� ��}���>�����{�S�ү��яcT�WD[0[������e|v��Z�!n��ۿ�"'�Gl�"�Nr�2���K��X���/Q�(Jݠ�gk�6�3�������V$pD��aK����Dz��yzg�|���������Y�[;+�xx�B��H.݄[�nkiv���S��fu�����媛P�SK$D��������
&�v!���9��|�J����W����s�2TȊ�+�Gf5:S��nY
g7nA���1�1&��7� ���Y�&wWbaK�t�6�K�ޘ�ch|��#���+�S�39�:!a�@���:�r�i��jm��lō���m�n�=��4U�=LZi��Q���T�;`<*B?q����R�}�-:4*)�����~j7y?�$k��P��?���
����F����~��)
\��ݓ��n^�3�nO���N��d�"%��4X�_�1�+3�t���\Ӑy��4YI��	 �,˭�"㻢0�2~1 m/���ѫg��
FؔW&x�����#"��K��i�WƵ9`�_@�l"�E�˶1ӟ#���]ӟe�%�7�ږ�Ɍ��O.�l):::���\�B Q<�w�j&66�GFF�~�x}�����9�i�,(�>�NO}����s��,���N�}Qw���4�N���ath���R����^^�H�WTăT��wC��E*n���xx��At��;��������'�~����#/�'35�M�B,uO	s�$,�\�	$�NU=�	�&���G�t�9�
���m�,�x����033��l��`�]g{Ȩ#� #�#��Kr{��+�7~� MI3�xE:�gx�9壶���[�:i���ؔo�:uzq���iii^~�щ	P~,
�7#7���-	��Q���v3sAh�&ԧI|.PӀEYY���|>�>��{� (5��D[��k٨?ը��.�ԋiF���+�#��A��h�m���
GE	j� Fx��kt^�B5��]/�y}�k�isWׇ	��h�w�Ts׷^��/S�ŀ=�ae�'�Whg����� ���c��lQ׏�[��==,Fv��T�`����J6�Kc���K���݄��N�V#FF1�ᑥn�G�B�ǂ�r�YY��C.��#�P}]���u�ˏ!ݕ�����EU'c�m�z9G�nW�⒒����ZVM Q!�M&(;�d����]s�o�l�fE����W�a��C��'L?��+�(������v��Q�4�`��v��H�&:!o�l��M�v"�|3���k�O�].}j�RN6����18�.+3�d��H���j�V��G�7�huy8#��ܻ*T�����G6����3E���gϤ��p�H%���$-��&+�j�ڀ���x���#���y#�%�?��xC��b؀6X�	QAz GG�K�<��6��:���)�����S	#Cu��Jpg�-����<��'�G�YU`d��=��2��7��O�4%ƺm�<6K�jB�l���/�_���DtA՝�& �uՀ�p��Ql��.Ѱ��if�`<qr�Y����$��t~�H}��p�*>�����G쳊��I�z��:�Pmb�W�HMᎱ1^s��w;3�h�K����"�=�'�K�L�h4H������)��ݕQ�L8fg���y�[�k�g�D'�^Tj�?ղ����L���d\70U�iޖpDe�wfH峨w���\��2�� ���	�)���ܲ܉�c[�f<d��"}�(Ɔ��������ف'�i[�A�Qd�vN�%1�*�\�m��_����s�|�u���#���V�.���T�+z"2m��)K}<�����$ڳ�iyU�oem]ZUն#�R�Q���o�M�/^C��3����;�_a�k������cD%k�lp�I��% ���1�-�}�Z�:ؼ��wF���431&�ߖ���2�a���w̕��FO��,�#�3��%"?�U��z�1А�k_e�:Qi�_��a%�<�1î����E��Ȥ'>�S����#��)���;`J��ъ|SEL=�<�#b��3���G�1D�!�l�����-�J�ٹ
����5&#�9��f�$j0q�S�d`���
uQ�<Ls�v��\:�z�IM�`�=��]���&�U�]t�������.���1xO=-��D+(k�)�1@��w������>Q�X���咱��9��Y82d���
R�c��k
Gcmǿ���]�{O�ţO(�{xY^׻���\���{�zM�G�f�ͷ'čx<o����!5�r�s5�W��D���ƹ,�C�� ������~���yi��%������&�#���]�� c"u���.p�Rm/6Nc7s�A�9>���e����"�+�h0�e�P��KMG6;,�V(���桉��_��[�A;���%��ݱ�*(��#��f\Q��V��b���"%�jz�/+��196�$ �#,���Q0^�&��X�|FĬ�m�����Es���\m���^)���0�4�5j��^'W	��p�����Ҝn�2S�ӓ�ܝF�����jf�4�c��-f�܏�b��Ę�D8c&�������{��:7d��} �I�J��k�*��3:j�&A`+S0h�l�d_��k����̸�e��}:�dU��{Q��7U��z��0��|;BD�w\R�#�,�4AAe�>�%u\A�/�G��⊫���^�j��CF���.��w&��_����6V�@`L9i�yBٓa���v�1e��#J]^i�[I��qe��7�+��X��P�:p��
��y���NyLD_�1&n�x5o�s�j�N&�
��i�0feuS�,3D�*o�ۡ#ѫJ� 	����w����]}��=i�?e�;�C���J���?�.�Z=���fyC�#$�%y��'B3�2�L��b1���t4�l��y���̌��������?�iM��\��}���c�����$�C���?t`��ҁq7��P^��^�*rr��>ئܛ�U'�����?|R��������i���?���9�s
��_��=](� �������
����ea7v�Y�]w|6�/PL��������0�_]��AQt�L�|�P�q�m:���!5^�d��x�L��@�!��%j���a�=A�i��l6�~��2/R*�2`�Z�����o���>��޺,-�,�7�8�Ms_�{Bv��&���vfZ=����a�L��2�V��Ӑ�G�5��׽������V�6����&��ZΤC��C�P���s
��K��k��,/�ʍV�@F�=�쮱�ZbLi<���k�����	��$�T=ti	��.�	菕ۇy�P��ا
�l����4}O�x��A�=�^���וO?)w��c.��l�٦+��?e��e�d��v*m���]��A�]��t��h#n�[�<��� <$�)'�\ç3=!%9~��J�ѕ�!�NP*��O["W�-�\���Vs�.=0s+ͅا��M���ҍ�ħ���P�9�W����v�5�ל��K�V+xw���_8]�\cg��]���b������̨�2S��%�$�?����w�O�%ٶ���1���2xbE/#.�� �͇�IA�y�����Xn�0�&)x	,���+��DLyJ���Ojx����%9y6�N���hld$�����ĩ��P�;�2�O���r��T�W�RI!����,Y$��	��"�M�2��-��Z�~Ь�4z]O���}fT�C����{k+��ZjCl��߽.�����+'�X�L����ӟ�0&ur����-��3~i���z|t�`75���mF��E#	vL��&��nx�~Qe ������J���g#�o�ߖ�Ѹz��Ż�.N_;B�($@!�S�6h
m���^v2�H�z�flb�^�Aޣ/m�d`�!;=3�3��NH��y��G��?��TUq�&����q��+W0dM���wXU��T	�b1I��d$�_�pt���E&�� ess����"X�d1��`b�K�̮��Xh����x��,��H��g 	�5���+F�/���3��_�*?�#ď�2Hs`�f�j'�5�d�x���g^ϴZ��m�+U��n.��Y�����~������,m� /�x��u��rl���]*I�k�x�@2� �Y������1IE���G�б���Q�g�{��T
��z�bH����u%{�'�Y�\��C)��[���Z++̿�l���?�&Z=q�Z���*灹RE����=��m8��F܋��o���'�z�51�4��y<��n�!�N�H�3<LH񖉘�_��8X���o�M���쫴~�&�p�&�G����X�{��)Q�AtN���'�it:1n5>2�8�:�
@º?��Ɓ�\���<��k��,���q���?U��u�HaR������	&��|HF&�ِBg=�w}'��`S��O��H�3	�[L/~����Ӱv������Sǩ�wb���˜�>b�sI�Fq�����-q@ʔ�#r��ۢ��g;�#��������*�ɱ��I*U�5�  Z�����4���Ky2|�?rث�t�����*�D@ 0;n�7΄I��H�Pzr2 ��p+(+?���{W���W�q*w�M���=v��TCբ��*���n߳�W�U��i(8�&3�6�ۇR�J�WS5{�l�=DI���\,W_���"e��?9&��kh�>�W�]���57��d���&�^ȨNN�F]_G'Xb�\:�?�Lś�w�y�A���W5����c��u�0[�=Z~u��=�@��8��O3 ��Z��_�h2���f2��|���]�jt���R�6��CY?�*-|�A��5�Km^ô1\��B�e�E-��#1n���.�tG��АӦA��	9V�T�c��ܞ�%�GKa$!��������f�� 1��Cw�4����@�T鹹ˀy�f����M:�
3 �V.��QO���b�K�*Csw�I�_Nbڽ�ԕ�J����?�ޢ'W8��螢���J�(�R��zt���^iA���]�<7C��il�����^m�=L0o��n���C�#�DҀ�C�[�������|���M��CE�s�nR��X���S�`����'(���|Gݓ@���IY��I�%>����=KP[��(R�tO��c=�
��аa��ቍ��������F:�~��(��7���j|��!;R�� �S�J�{��=,� �"!��ZO?����gg��Ub�&lA�	ޗ|��
��9ϯE�$+$�o�Q��G-l�/t�&V�}����[�K��RL���+�<J\Tb��_T~8P:��k�I!@�6�jt3����	d�����h���GEE\��Ry��O�K��X��}��}��Vc�U�&�3r+n�[�/�~f:Q����� �A��.[�}���-G�#��m��h�`��GR�T�i���l�� ���TR===yƇ��H�I� \\���8\'�n��ŗ���(�����N�R�5mB�����#�;,q�����%�D��|~�3�u��E�6S���>E�l?����_6�r��~1�=�>f�;���@>��ʊ��<�2/���:���i[�FJ�P��q�O��f@�a����E�:�V+���?yd	H\��w,q���!�Ɩ�źn*Zń;b�Ն�/�^.==������t �s���J���k��|��M���K�xG�3n�?(f�����Y�\��;�v�87��cC�V7����?"��e�;#'���rtƻ�氋l��+P.�ouA#��NOO���Z�Ew�e�9ύ�����T��&;���g�K�$~^}�h}��/���a�1�������ݨ5zg�k��)�n��-?�����C��8 �L>#C���8��>�n�e��ݘ��M�j~k�xza���v��o2�2��(�[�Ӣ�D<�OtRe��_��#�G�o�4L.�N\P�]���}�-�{}��a:�I[[o�z�~/S���vtt|h���b��-�4�4�ý[9���<�~_T�YFd���o��xE�����Z�d��yS�o������S�f��w���%l�����������3C���ꬡ����ï|�zW!3y({{{9P���kk���Ñ��(�p���x��U�%�d��;��ώ��������2*�1VҢ�n�b<&�F�����0�������� O�=�?-r�؁��K���r+�Ֆ�������;W�y�|҆a��uZ0��đ]RP@{M��v���v~3��>pWr�9���F}�צb����}A|��omm����"�IL�^�>��y
H��iw5�̤��ښ����*ō�\��<:�o_������SPP^{L��j�F;����;}
6=ݷ֟���[R���F�.���{�7�������-�ߪ@��]�^=����ڂ��A����j�Nr��~�z��B������|�a������Ω:kxs.i̪;س�����.��izy�m[�9A��n��k��*0�ߨqA;��e����<;Ȁ1�;J�W-�йrħ]�gU�|�]�P��В�1� �\���v�����v/wz�8���e#�b��&����ރ�d��$�r�g@9�m�@y��jJ����?Wq�>���>���e�t膮���u�� Q����q8������,Ⱦ�ݫ���yxvz��=O���ϕ;L�R�����zg1�i�\Ʀ$��~R4-����G�>�� ����E$Mc�u�?��d���"�&IFEA�_���ܒt$>���?:::I)���Y��"h�@kW~|��bsaaX�k��m���Jv�\�8�e�4~�A9W����"�o���-y�E&���N��W٢��5#���=.)��H<,~�ɞ�@%����~��ﮘy[��j6�.z�"�쫍��$��g���w��-���z��^�`o.y�&�.\>�ذ^��Ewt$�~�b�>VX�כּ(�a=tJ�������4\>�rH-.f�C�_!��$�u�*i�jd؎D`���'�+�fzA	��W���"�}2�.���R���UF2ȅ6��oQ^&��ej}��v��۴�Q�
k%���lk�x��Z8�'��S�I�QTU���x�?�ǟ�}Э3���f����>s���!�+

�ۇ��4�F஝����S�-O��a�xrm:��Ϝ-�~,�O�0'Ǻ��_kCн^8����:�]����4/�O�h�}���*�7:�dFYE�8�* � �0�A�)�7�w��\`+a��ĺXPe��4\>x�>*3�~�n�~�H�'�I߭�{��&o<���Y�rS�f�P<���W�~�J�2�ܚFJ��$�� 	�)����BPP�z�Ŏ�[c��_	&�A� �E�]������4GLQQ1f�\����ZF�1��[<7��@���2��}/A�w�0�4���}�吃lJ�����#��Z��5�����u��`�?����	�:=6� �MJ$3�x4|��Sӻ�|pQщ1pL��!�
��_%�@�Ȭ	��=���{��*z�����n�D<`�3�P�����\qm��:�4O0%��(��찷:Ǹ�:���kK�e�D�w>¿�2>٭�o�]�}������#���������`�i�h�"�7!����'����#���(�m��i�%�_����;UrDu�����Z�v�m~SM�����nx;��;�T��ƈI�t]�~b��0�u
�G&�dF��w��.����@�NO�	Ԕ���}M\��2x�˶s��kkÏo��+U����7Of�w�e6�v��P�	� �dյccf|퇷�T�8��-p��ybBެ�KU�#X�e̪Q�k���B����T��sj�pq� �!P����.1�����r��А����`{�{$���s�.�J�^6߬/r�XƸ�)��"�[��r�������VN�XXXxs�����*��0O�5I�(='���'=K��+��Q?26�5��T;��2u� yDhS�x ��7=djW�Q"�
��}�g��i�/����d����"��uHn!�a������D$���z�?�L�[m�u��Uj3G������t���#��pКBs���ݭ��-f2��ދf8������?C}��-��vj�W�n��e�������������ܛ0ڛ����ڞ靏��<k3%�g��Ǉa���b��ink�b�h�)�o��6EZ�P�](|��������Wa����yy�
\ٿ��TXX�4��L���en�[	��M�N�j�2O#e�d�T��Nr��`kD>$#t�V�إ�r���02�^�B ��M�#ĭOF�%��x���-{;���]ub�2!�6���� T�G�nTZ���? Јhy!��8r�n�Z�FN�h�����
qΌ�ENU�76`#q^�o�9.�H&�t�S�2�]�[R�zY.���Y��q0̪����E��eWF�F��-R�B����di,0ފ2�
'�訔�4���;��h�	GP��<�"V���[��޽/�k�[Dd���o�I
g�W�
���C+N(�[ �`��2ppRY�=Н��'
�� �@��'�����*����|���7��nTx�f���� ��Z�"�F��1>dj�U�2�9�oi[������ǁ'm�`ü;D�x���l�r�����Я��ąߡ˵��SAip�/�ܮ���Yvcv� ��<�����:�X�15���Wu]�T'�y�ů�͛FNq��A�_�c;��*)�L�8c��<�q�Xg�GB\���"OtA^�����l�`iyyaee|x8&����D���mjș�B���y�c2�#�P���a@��~��c�.�UϺ}/���`@먂���ek���͑q��L{IJ�f�9��%�cEL�'l|�I��O�H�K|+)G9���3C2���7H�	��8'��(�O��WS3�.�n���ge� ͥ�Kg14S� 9  �Y�+��z5h�/�sT�С�;f����������n6I
FRCE\���+�bnf�~�������w�li��׎$lhܯ؍[�n#"#?�4V*K_�i��]��OZV����h#go.��:�)������ 煉����Q�ɛgT����*u��.ȿ�%��>ɗ����l�=���/��a����s�k�9���l�Hl.�T�F'��r8�N�ACC�9eYޙ�jp���W�L��-?��^D�cw�˻XX|�
��	X�\xA��@��קTVV�$����e.��;:;1noo-�,�[��
����qh��е-*.u�i��$�[�T̟b�Ϥ�.�QRVq��Z�@����������R�L�}���ab��U�3�Ӏ��x� �[��aC=�r�vtG����NDv���4r��/>4���7.+-z�!w�>H�j�όj�K���p/�����d�|�TV�@"$'+���9�����X����{\'ƛ�d�=���� �"08C�Y��B�y���l ���E�!Kr��Ѳ�Qs��Ӧ?�����c�{Ł�����>66r�M��w̮n��x'=7�5Qԗ�=����0
c8��0�#.�:wP<	���!ް�.~k�}w$�賄�+q�|'z������K:;��KeI/<כ?¿�i���t���4SIIɡ\���3-���b?����� �F��kJo����WU����*Ø�m�8>�i����p%����&+˷b|���;��Ld����:+ַ�1�x������Rf5CLh��Ѫ�r�
���EM*�����
���n8�U��1`��~*w��e����=W�h�����r��������g�SA����*L��O���j��F9V��-b�󵍃�>N�������u�Ҭ�<�`�^3�����h ��t$����w�x�҇����Цc�F<=S~?+��G\�2-�� ���݁���Lܪ`>0�B�]��'߹u!^#c���iɣ����K.2�c�O�;�YsoY�p��%��0�e�zUDNMmt��b��U܀�kꝷSlk��U^Ϛ��!����u�.����Ϸw�c׈��$��w��u=�W^���@Y{p��[�c���i/�?�bĂ�a�u�TIq�̲��o������NEa���=ʖH�{�FB\�-�sp�]���������e���a����إ�w�uj�D��!�ɧ���0��YE1��<FtQ�%ʾ�A�?�Y�B���(�.��Z��L>Y�]o`O�����4?�"$^2�i8�R������$�u'=�p�~.��S�,ꉀS�*����e������5�G,,32��� D��eq��LOP^$�*9��.l �r�\��y�%����!~��"��~�5N���MS����ٟ�����+2R`�z�g����x̳g����^$G�L��ʼ�)�!���~�Z\���R��X}��9*B�)p���9�B���
�Z�yɜu����3e%55�C��7����Nۜ?�D���x{�d�v�oJHY�����J��紗.$�����|a#B�����[$���q#Hy1��.�|_Rq�|q뭚��qQ���� ,E/b����*;��+�����*��Y��))��~���[���^[a��i���糼N{�5�35��I|x��f��T_��Y�"z��")�[�u-���"G�r�"0�l%�bwm�����������B}c��f��R�H������3���W��C���ߑ�80ޚ�Y�s���\�C�������¼���� I�"�[��|�T�<m|ˠ�N�>d����QK�mo.�YI��-*����.]��ƓM飢Y.�7��/�#顉�r��&�������A�����j�u
�j㳊"��&����b�,#�����+�Pn��+�c���F������ �ն{o;����m�x_Ѷ�J�*�ϴ/����)��d�$E��\�~��]� K�IM��mBD��Ě�%>-���$U5���VM�pB�]�lall,'??��	�W���v������sݹ����T3 u��9���niCa}}�	�6W�\�} #��|G\�l�(K���B��$��]�E����m�6s����f�Ns�X$_���ն��Y������u�S����������P�6:�q�j�@�O9�b�>l]�l�x�_IEeH���S��վǊ=+p���WW�!1�h��7n�X�u��
8�o�&J[d.�C��S�@kN�/�o&�]�:W#س��y�m��oD��'qd�"���ތ�U�;���\�Z�G��C�wk<�3m��|��j�vo�޽��EP��������,ѲG��|�X���x����4�mQKa>�ֹ�_Xm���T\&��KV�������~��j���w�H�V���� �a	,
��/�A(P@���r�|�^y�#_{W�~>�֟4-�M�Tn
&�.��^heP���;eB),\��X-{zj7:=�7w�уo��(}/'.u�X(Y�&� 9�|7Ⰻ�n�.u<��;�9|�]���#{�=���o����	���D�=I$	)�f��4�sv�n�&%@�@3�����n?dffNxH68T;PzQ�Q�ѧ(���G �N�ݞ��}�����R~~����c-���bؚ٦]V�e��,�3`;3����o��W�$
���777'���9�+���j�0O�@'5���1��4��h�.'�ZH�������"���r��j�����]-��r�w�t����-$PC��Ƨ-�43��=���ʻ�dViQ]Q�T�6/M��Ν��tC<y���}��*�:n%�5������rrrH��,j�y���5?ν"z$JC������TIuM	�<��F��9J��X�Dv�&���ョJyU��<n��9eե�=��^;��67��5>4��aR 3�������9�#������a��:�M�v����&�$܈�hڞez� ���={���A�=�l/�O�G�,�:�=�	��15�ʭ��\L�I�{�!�B��4MJ��0%�Tց'���Q%�P�4��-�7[0t�TaΔ���&^	w^��>7�Yx�V�Ǫ���o����Ē6�Ð
��G˘�LT�Ő�9E��U{�]�����L��g�R�Wl<�O5��W"�Rۛ�D��o-6T.��tlyP�d�S�c?�=݂�LX����π�>+�ޓ�����_�P�x? eHi9�t�/�5�&�{�P�5���>���֮���l��0���F;��ȝѹ��?+���SnE|;Z�X'"�-��tݎԩc�0)͎�.���:�����2���	}��
i��_HE�y����tW���~�7�,�Q����Q�W�'�Zi&l���#?w�2�
*ͱ�\ҧ�����u����b����9�mN��5���=/���2���9b�������,�SSTՉ�",���z�Gi��lH����-�4��~���S_���*��J7��tI�J" �%ݰ�����tw/R�,��ݱt-���_������y�p�ݹw�{�Qc9�9h71s�m^O7��y82=!/��؟����q��`�c�O��W�Š	Q����MO"o���m��;F�,�����TUU=�����o�b
�y{����f��ٿ���ohh��UJ�c=��/F`y��z��p��B���N5*;㷛�SPP��1J�;;����0O�Sr�V�
%*�Ϸ8�::Ze��w4X����	WG�o�v��}��!�:�{�����Aw>ˣM��GU�M߯���V��y�F,vJt!a��5��`q�C&���\������	���1e?��ԙO@`�壛J�]K 6	)E��P�v­�!F��j/J EE444�������L7�_����-jV�n�c�===���_�g ��N���E�2��ٷQu�m�(ǋ{�Ŋ��;AkV#D6����9��nB�y��� ƃK:s�~9�xkS�gX�*�(2�R�9�S���F�GI#;�W5���u�ܤ�?_���[���q�&��.a�a}�o��>I�e�Z���t���;Z���}�|o,���N���-|�O�i�mL�fM�e��G��F�~$�2�a��:�����r��&e㤍�t�� g����E�'K�ZE����j��O��7����17�`0�E>�Qޝ
+Z�|a���^����11b/���}�"�Rs�_w�G�	fU�I���'�__���p�{�J��~�ߨw�6���0uP=	o:�Z5@�/x���>+E�ݞ6� ���{`wS5�/`΃Q��pȂ�!��@Zn;x��-_G�g��m1_*��ܧb�mz2�_���B�A}E�~�j�fpdq}�@��܅�@jSW�>G```����	ؚh��}��R>Mi�T�1ޥ�@�e/��/��s_����=�Z��:Υ:ރ��H�$��{My(Ž�n���'çgO����3��U8_�^!�^��7��u���}�t�H3���\�6Q���3h�:h/�$p�?�Z�<�\1�8ۭ�E6cnz�i�x�� �<�2�7��II������:,5`׶�4�+�'at������Dd�Z5,L?\]���� |U�񣼜{ %qI��HO	�J��N�ce�C�$Q�d7�og%G�r68w��d���R�^lMS���\�}A�1��(�1�	����թHb���yc��8<��n�Bv�S>-5>�B�z�EL}�K5u���a�.���yZC�#�SO	�C��o�
�o��7<�|�LL8`�;�/���fr�+/՟�}�Z�Z��_�L-w��CH�j������� ��m;u��08�&&zs2��!b��#�%���� ��B��(�M=�D�d7��w�v�7+`���,EW��<zEj^I)�?	x�#���j�n�X�������X�>("�&{抯A7��.������r�3��E_f��n�#s���j�]�A�|$�b>��:߯�3�u�Mp����@b�T��U6+�B���]f�[;e��'�p� mǽqtXz=���%HM�v9�f���S���uzMUy�o	}���g?�}?51�I3_���r��a��-Ob��pYyyT�o��K6�'$(A����"�&c�fmA}��9��ʿth�c5���<�8��Gcb��M[Tܓ�Cm}����$�������a�dA�M)㷧Y������z�v��G�T�����5q�z����7Ř�*����4Mx\W75~�g�������6�~H:�����[م�D�x5荶��M��0);_:�0&��̶�;�̼{����ޤ���\�����^t���^}�E�뎋�q��AW�PD�$sG֋�}����o�[gӥ��MLxq�MLw��<D�9__�l��۽�|��g��~h1�bb�����p�
Z}��ʲ�/��������;�q�-����G"vvg�C�K�����LZt��!��,��2�u��۟��qf5��[ì�KG�322�a����у�&?���/~{c��.w��x!_ǩ,>�����fK7k�V;�hh,f��M�A��l�W-`[r��5�p���G��݇T�_���eڿN!��*�IO�	����O����l�~~7�>Q1Z)�@��u���vfvvk_�Й1�]�]�GH^&�{jzwwd�8����dº��oF���"!)��iBI��������y���4%���h�xx��<Q6�iN,=LJA�D^n�,�+�G<���tKH#���͚�1N��	�������ڟ,`�q���kK��r�F5�k2�:99q�<^���+k@>��?yo1�L��v`K7YuG4��fN�IRFv�u�S�dË8ezM߇��`�L��UA ���2|�69�Bvx�	mH��Cq������ ��W�e��s^$�eA--o:::��,	JKK��F��fY���׺�)��1�47�a&�y�/�tЕ�,��m���F�{o>%ɜ*�.ڴ��j��0�r�����'m#^��-�a���w�f��<LG��@�gۘw3Q!���z0�>]�����TF���x��HHÞm�����л�(zss�Y۸YPc���}���325��!��\��{ra�|s�U�B�*5���x}$�}�+'^�ׅ}�[���l�r@�g�#Cе��W�������9^� u�g`�:(�7A���~+𼺺:����ejn���h8��d�]7k�|m���Y�w�������och[��hx�B�i�#����~�>U	e��z�RL�����!DxAB~HQ�#��.l�z$�(�k�-�i9���2F�.8��~�����s��Q;�t�!;�M����`D!�].]�}.g�̱�5�A�w	>�d�Q��+"�=����X�e�-�����e�<ݚ_ڕ��ɧ�ƥYb7�/�u�M�����㪍�Y��)�wƊ��,����Tk4v������N��@ 3��BB�(`JJN��ccx�E��`�#��t��VV��b0���x�iBw��y���Vt=�*r�v�ww���)�_O�I���V&�����a�-##CJI�BU�u:+I-y:V��T^:_o���
�����5�~���j���h�'+C=٫]hH�/������(�����������3��I�E����y��qö�*w�SJ����G[&J��H���6?���	��\��ZZ�9�V�h.b�q0?w��Zv�wrFm|J���ʪ����ӣbgg��珛��#��674\�M�.Ti��x�:�L�V��tnoىHC� cW! ��k��,����`b�l��N��S?� ��X*[EFV괎�V�e]���f�����Zű��M�b�v�Q��/x��ō��J擳��nS�T�(��� ^�}��{u�Y07 F�Q�.�y�"��Pp�z-��E0���]u���}g?�������F�ދ\��(�ޕ��^<�7����s�i�c� ��k_�z�|�wcS2��O�DK����˃[�����VMUt���Q�e�A�͈��]�ZaX��J�	�kq�n�D����fj( �TS�C:�1�������<�k�U�N��!H6����Ԥ�ݤa**�Q>�:'�-�/���9��(M�[��张6m��k��=oHd1�Z�/g��'���3�6nv�$��@�å�O�B�Xg��|���M����7���u�Eo�ģݿi�^:��b��+��+SfVVƀ���f� �P��\Β�I���xK�3l�R?	L��|cGh�\�{F*���K	{mIL����x]b^/5t�%ʝG��>j�ч~8�WA�S�r�Y�2z�ɣ�d����h�������H㏇i��	yݦ��m�ͫGD��\8�e̜UH���Σg��5c�]]�ß�P�f�X��Ƞ��۱�g�v��a/��@C���h�",��� ��eRXx8���杺: �}�0ic�ߒW�zpw0{��bЀ>�'����q� �Z��7��+�j%�!Yl�7p��T}�%��"n"
}l�~��;�$2��#�~$��VVƝ#���O�S�a��y�) Ɔ?4�r�6���4���ַ��'���8$-�����	0�ؤT}���z�ڥ��Ы����_��g�I��IQ�j�G��F=�3��ON����肨U	�u�͹����=f��=<�p)JAϖy%e 7g	k���o�9AQin^^�I����B����+L�N骋(�a��eJ���v��'"W�[����f�tE�~/Q�A�~�l�|�}�m�8�&��R&����,�=?�`h��nd) 6�
�����%f�\��}�&�(L`p�)�l���?��Ǧ�X���������G&��	[�ӊX�Yx8A�Ae�4��oUq�w���]�\�����a�j�`��4@���������[	 ,җ/���7R\;<9Gx����(����B����v 3�Z�0g�F��'s�Kc1�
���#��b�%���8qڏ�TQ{K%@�]�h#ܲ6�Ł�����	��:#��)�1y��xR�)s��(�Qw������������+˵Ļnd�+��8�[a�F�ﺑ8zK�ȑ���t $�d,�w=��A��������䙂�&�p��gH��&o�=�$+,���d�kEE�U����(u=5g��夊) ١�7�#����0xJVLp}�C��+(�=K�}=�ؐ�B�ơ�K�LU1}��{� Y���e��$3����-��� q��!��{ɚ������q�>�jZ�tIU]	ŋ�>�Cd�}�'�}�iJqm�-t_�hE��^�r��|��B�0�%v�j�P(�o%���e.�dm�]dؼ.$���kÒP�X���2�Ϩ�麷BQ�\�<Q�hУ-�Rd�R.�(-~0W�Z�I(��+ە��c, �A3A��Q����i']]�{�ZĂ�㱚Ǖcx�%A��#9ug�肆?�Ρ��Qp���}9�+`�ރwooolrr���BY���&�
6ԑ�(�54��Pn$�n'��eH`�jP/}jH�;�ns��ꊧ�`y3���a�iϮ�S����nݏ-8Ӵ�(�Nk�Y�p]&Y��1O���kd����f�炋�X��zs[��<���g��\ѣ�6�\ެB�#^�Mk�#!%��nmyU��i��ٛ�[���e�����"��lD3� ����r�6���iS�c���	4��K 3U]��4=0��/���g���D�*���S�0��_]��U�oٸ�z6d.��u׭��$�n�����[̺�CA�ۼkvb�F�c^���H�RB���[��4��ĥ�|i��A�>�q��Ik��Δ�fR�
�w���&��-��{B�F�_�ʀH4�#�ǫ�J�ɷc�����2F��uK1�>a��ec=�-�b>�_1��de>L��(|X�/3I�E��'��V���J���7}���!��C�T�q�K�4ES�&e��m��m��w�r�&�#�j��b�����^��L�W�c���a�����1"*E�E{R*����ǚ/�(����d������D9��yfU�+�w����f5�&x[B���ZM�5�ٝ���������v��,�O3�
ۄZ���jZ��ѯ� i^�����\\~
<��*;�����-����r����W��M�%��V�Z:u/�i�T<�?�6���y�z��Ҽg䬥�4�����E�?���H"�;�T앲,21��5�R�Ew|�)@�x3�E+�[
��4g�ᐴ�#���l�vL��|��X\�y�mO�.����従{�qM)���瑢7�K�Go��
�3�:�>�K��Z�[����@j�5��4���z���pg}����$O^ԉ���a__��*��9����e�}.d�;���9��y)1��������a�Q���"����x�������j)�i7F�0��{7O�����[��D�/6%��~K�@�T��y����Ulj�.N�N?-(FK����-9��p^`�����5��#�kR�+��H�4ة�
�}+��g�Mz������W~�l��k����eT7�u�����5Ia�YI��+����:�����#��ĪI���D��+�G�Wcx�i�M�O��V֚�o�d�����@���f����^���������G�����������Y,��%$��D��(4Z�WRf!޻��@̈R�a�7h}r�N�+xG�(G��|jf������>ta'�Yg5�܀���!���C���ŏ��&}1�$���d1��	�ͰU sU��C՗vz_�YW*!��zr�c�:L�q7�e�Q����旱f�r�cܯ]�S��\��y�6�'O%��_�������I���L%f;�aL̅F�w�{���s�1������ZLr�o۞{5ԟ__��-,>D�]��P~�f�/����ik�u�ϯ��@"N{���\պ^wD�(IN�>ǳؿ��w]D�G�S�b�8}��9��(���c���G�/f U���ۚ͏*;�� �ۅ���VS˛r_�Ύ���ۉS�3��
�{�����u,��L��M�Ln�b�Z���d>0���2J6��NR�����x%�u�<(�� Kс�#�MO��99B��.�Z#�\��.�-uK�q�����.�oF	߿V!l6�Y	)�*(� 	;qx����Hʠf��q�[O���0+�-����&4�O�6�����<׉�C�$~oP?`��B�?yX],�=^�0*d�����d�&�gm#t� Ƣ��XIE�.��m�E�7�s�=���ᏰҢ>��\�7�lrI�ۉ*����g3n�Rv���G�1wXJrh��G!0��6]�t�6�@m�l�QdU`!b �0��StJS���HM��5�Ӯ;��ҩ�����rSS�c��}�N�o�q���\d�
X
M:�"�}TDb�zX�$�y��T�Ww�⪇
��q���
���Ռ�S�ʷO��$\�N�5�4�����J@�,���G�	]8���k=��Z����eo�[���"����o_���p6����[Z�9S�H?��tO�B��酓�H�����G�:	��=^��!���v�U��vi�q�HW�����L��Rsa̬;���/�p
NP���~7�e��7,�)�q?�x3f	�z��/B�k�&�������i�D�7(_�Ȟ:��K/���st�<�S�L?X.��)�������>E��e�ѐL/ה��q �[�4�і�}Op�4Y�n77%��m9�QZc��Q�*kQWm"��j��#cr�a~�4ߖ����S�>�n��}k���Ͷ��bҌ����Ds%��%I��_h�I�5��0�Dm��@=r�NR���G�
������ʥ�j�IW#<u�΍-*��&Zµj!YkA�E,�&&8xxY;�ԑ��Am��[3`�Q�.�`X����bn�~|`]�
��%�۞�KR��D��kgI�~���o���7	1�UPy�'��XV��cP��G.�����x`3!W�x�ϝz����zҍ�	�
��'�g����0LW�;��
����J�3��4�Jh�I�#	&�u��!2���΂���J�;��#�� �U63�xY<ṽ����f���B�yo�a�d�Fr��:�՜p-X�
ܯy�"3P�Z���#|��V/2�%Z��W	�*F��d��j��
Rj��]��߇��|��{���c�U��|.Ð~y@��W7�,ԃ�d� Yu����"�XQ �v�- W�ƚ��=����Sw>|�J#H���ι���A�����h� �Q�?	��K��2���Wqd;燫�&��x����H��u��9px�"����0�@�q��ґ��i���ݸ�p��	�ײ^"���5ɏdk���,GFF��T�W�y��W�����I��:쒉r|M���5'x5������f�n�N�#0jn���l�D#�� X��,x�5u"�|F[G�1&E��;�⓭	���bt���v�����9t�tx��e����[����xlE/�9��0%�K�z��Qg����5dԲ��B:P�jzZ��
�g:���G#�q��8/k�P��gSR�ߦyx^O�5���KV6�f	#�2�P�e�hɩN�QF8uc�9�`�V��^�8�
AFM&=���V��Dt��+�J䯟P�!**w�������l��դ'����μ�e$�X�݆Zĵ �W��cY5P"�T�lwF�1f�kxR>2M� B3�x�I�dd�z�`�>�_["�;7��sIIoO�T(�%.����r1��{��D�hq=�����\o(��}x�/�ÛCZ�rc�h�f���|�9].O�o_�\�?��g@�����PZ�ۡl������/&���&��}ow����7ww�	�2����)���t3�����e9����	љ����46x}WTr:)=0,��Ti���*����=G�c��ŀ��"Ʊ5���O�z��tJ(�=i(�����؉���\��Xp�IT�ggݏ���6#/o��^���)�ѥ:�r�P�ފ��O��%���7�U�9ά�s�~�������"<�::�q�:���$���"jk���+����'x� ۻ�X=L���p(Y|"4��l����ׯ�0���k�G{}��A�C8ˇޅ��������Ԩ���M�#i���J��%�bAʻλ���
v�{�-�4L>���$�g}���R�TZ!o[=��s!���L��e.UUUz��|��e�%�:�G�As�R�vK�-N��N`����-¾��c��`�q�岁*��h��9���J�*0����p<kw7�s4_�$���n�
'!�Svt�gʫ���_9�_�D�ӳ�V����HD�E�e5�}}K �)u ��V���'qMKr BY�4��Z��-�)n:����z�m��G+��:E��<�~+�Ư�b�n���8n�ӽ�$�� QѼe(J�߲�b�� )�l%�T}��t�g�l�ʘsѝ\�g
.nUCsch��?5��E/!o�SRr� ��]A�ZW�V2��	�Ą�����ͅ� �C,%��&�7B��<Do&SS��2�����Й�&�.Q_P��!@��JS{�8s�+ό]5�̉�����}��e�]�����D��z3��p�}�r�R�}7~	�� QNgQ)
�o��"�T/h�KLOf�������NOI��2�6qq�n�i�.�=��}r9?[c���K���6���^9��S ��de������^U�z��So����7�p"z�>��>t۟�.Qﱶ�:��BQ�q7��������ms��B��ɑ
N����ͮt�d����G�G��h&S�s �z0��ЫF�li�-�	�1j���N�zd��u�o���v�tl�H��R�_V~�Ȕa���w�M��R�pԌ>!��ymz#=8��Tlכ�s���nv*�E��� �濥��(]�[hHY�D�()=���x���0�_a�Ga�8�u0ג���}al?���LL9P&&��O���c-�\��l�7g�&�������肬�3Zii��BC۲w`�������Ɩ�+�a���W�)��`iQ��$��h�:15��3�rV:uB�ivY�,�~}��y��b�_��d�Ʀ�j��@��MMG^�ލ�#֜�a��i�-l��[Ǝ��aGi^r����^Ü�g���O�_D.�x��^~�XjE�H5"]���'�cn�uE>�,^~��x3U7!�Cݞ�᭜W�]e���l7Js���$��/ٲ��H��w��,�:�W_Ckp�$}`�K~���\5����~�tF�0���̻���N��Lk\��s�
_�L��Y<�{��,��&���^��iFZ/�	IF,�<���\.�9і�.���~�w�$,�4�GOիj�����9�2�&����������)���6�� �1�����mmˉ��[��FK]��7C��)�NG�i1�o{�L��D/E��$\(�ڿb��Ku��jk��'�����2�\c���N3¿�El/D��-��I/H4�� ��)�\�*`�GJa)}�L�	��	�w���y�r�������~{��j"C�[�"�PA��b����}��_�d�~�!�[�������m�{��&�C_Q��iy�����ΐH_<jQM5����N�[��F�n"�Z-��/0hW�Q�`r�?����R�m��+A���<p�ޤr�>Q����6<�o�O��>�|�����$�-�3�x �F�0X��9�� ��7@q�{��CS�q_�.ԑL����no�*��'��g��;�1{'))����.;	��Ү��`J��_��hn_di�/�9�"H~�Y��u�F���!=vY�/bY�j2y˖�x/����6�������#�]��r��G���1��m�MQ	�;�a.������R�8�k�Q���5�\=}�������,kx�������&�6'�;bo|7�Sa���z�ٙ��U�y���(^I��Pd�iL��%��s��8��l���X)���E����B�K�⣼j��ɂ�@�s��*KU�R�AYB~ۙ��H�.]߮����J�'�����x�m8�B4z.e��<��z4ϕߏy�Ez�Д��_�]�'����!�E�۞�`&���?���g���x貈I3�l��N2�2�Ic�;�T�&�����j��a�M�e�+Qq�>}$��#���ޢ>��-�)�F�tF�m(6e�:{��4:F�4h�a9��2G������cKh~����{�:
N�,N���	Al������\>�4y������s1��`�n�xP����3B�'d�9��ޘPw?ס�%�������,��0�'��^/Д�cjkk�w'*
��:�g���RM;`�1/��e�;{�؟��l҆�"�x�O�Τ��YQ+P�^�7J]t3�g�����#�m�.��n.w�0�]�3���/{Kn��G��4!iهuE+P��0����<��/4�+�͇��Q���:�t����J��d�h��C��s�����cS�)�f��q�6m�&��p�!�+nq]k�@t����!������2��o�E�l	/�Lqq��WݪҔ�tC-]��	�۫��N�3��o�a�fr=^;9��c-�5R�n����r���n4���Tk�t��=��������|����ϕ�<V��G�π�MR��E���R)�b�%q��a'��瀿�]����j����j&��V��I<I�ԇ�O.�B��0�ۧ�V�5�ۮ;,��.�eS؜k�P�
������7J��2��
.�@(���-��<{����}aC��v�|�H]�=	V���EYE�G=Q$I���K�SD��,���L����K^4�+-��l=!MeŽ��$}j�D�
aJ���]��# W�3����}���ར����ER4�h��@3�z�qK��hIn�Db%�ihB��������ZF���K)����77Pw�ډ�e��dmG��9;  ��q���͘2�S����HG,�ܞ�;�-�uB�-x�0e�w,Q�� �޸���!q%Į�
g��5�&��bl,�Z� aO/6�z������Fg	bھ�@FP]!5젶/�[���TPB���Ƥ�}�m9�2�/?��ٓl�N=`!�M��"W�g�,&&�K���Q2�?�H~�%��7��>�1P��l�XR��mB�,:a>�ѿF>;S4X<��z�R8��B}�����{�~]�ײ��jj�L�7���$�I0��)��;� �ȏ��;�<�J� �l�]���1�C�܎�Z����i糜�SX�E�z3���-�[}��L� (�3tq�J����tTZ�-_���[��ϖOe٪��ڙ��WH���=��pSFl��+Y�Ϗ�N�9;S|d�q�;��Z����_D�ʹ���|�-_��_�L��	C��ǣE��C��dف�'B70P��X�x��[�f�n��yPv�x��W^���������ŦO:�DC0�޸�Ų�1C����}���}����*�s4���樔�:34|"�_�=��jqf�Ή�3H������ ��a�c�=k�;h�P٭0W�MR��e5�l���c��)	p��i�ܠOJRrFhe���ңm�3=���
S�N�eX�kBe{P���W"X�o7e��=.ޜ��������"8��<s�øvT>����n謡'\�Am�Ń�_6Rߎ��j�x�&�1!�~2�,J29{خ]�b�?�\��޹��(a/�_e�� �ߵ�$����X�oG%~���X���G�Eϑ7(1f����M�3J���i"�V�2�����dŁ��	e�H^t��~�2���.��'t�����Ϻ���Fk�>�v!�@��x����Q� K}�p�WŮ�,���RU��<��ON������1�`�5x��B��::H,3�O�Oc�.B��H\�37�(?~q=�h�z�R|d����<h���c�A��w&��s���"�?j��P����᱂O�y j���}�Յ�Χ���IsM~3���w�)u?l)��j�w���q_����{��fz$q$��5��悺C�z����wN�O��6�D�+��,�A�N�K��zĦ������V���D�AM#��A�]�EL�gOB��Y�9����"�3��d�e�,��Q)>=|Z�_~7����ݲ3�Ť��պ�>h��*B2�e�����K:�F�{68Aе��c�J�Y97�����F�!���c�֏�U�Rg��P��?R,pa�s�(ox��Μ�FJ]�~	d@�Y����? 1uņr�B���H�ݻ�dWc���^Y��������f�	r�N�ϫ��M�5��R���9۟�99edbr��~TܹJK��촞��Q3YwO��?]	~$��Z�a+��Yv m]��%�eo�=h懝&1��;XIq	��N�;����R��|q����u��x�ry�D�|D]W,3���#��8h�u��ן�����k�4�3�����I!?[��c���UxK@@pq�üc8��ᬁ�7�
�΁��Iդ�jXe�\���P}�?��P7nn����zzzÓ���ȣ��]]�E�یF����vHeYI"��)w~?@�SZ��5����F����D���_�7``�L���yo�^�x?]�N��z}am���s�R.�[RSY���3f�>�(��M��D�"��sJ~]�"޶lhcf;����	��B?������Uk��jM%��Y��K%�Ɲ��G���s���:� ��d(��_h��D�?R]ĝ3������� &�&Ѳ��{~�ȣ콿*<}=X�㳭:'2�=�YG-�k�CN%�J��@
^���{u;�yc[[Nd���)�*�����p���w��Hd��OQ���׫6�6���m�
��"< N��@ �v����-Y�R$���f����>����,SK'�Ș�vŽ֎��%(m���LC�����SҠM�zeӨB�'�[=�Hޓj��R|M\��
M�"����K�G�e
�{�L���m���>�t���Vչ�H��m'8v�g�+�$�E�������ⳛ��_�rZ��b��s	
ְ��KvT��u]��w�@W��6ŏ�m�U����Jx>n>�O©��9u�*Nu�&��0�K^�����?�`b���}�Ko���Ə��tX�ļ���l$�*�}m�J^	����N��F�/��������ڃ���2,8�7yӍ6��H� ��4��C�4�������ӌ�9o�r�cZ*�Ƭ��)�m4��s1d�Ϫ@������]%�CByyy4V�϶��G���h��X��})��g�Q�?�g���k��ޔ(��O�ע"�VA��zQf_��/­��~�+
����A�|�/��Q;PW6@^��Z.��i�;fX?��Rα��9���}�}RU=|;e�;͇��4�l�7|_`!c�n�	BJY`F�9���.�	1�B����i�x, /w������G4��yGG�1��y��O��o4a�$�4��m�)�	}J�Hߕ����R"�5�B�rz^uu��AS�����`{g��[PRT$H��r�w�P����ƫ}�[�MB�b���m���?����~��Qqgd�jRj\����A��q���W�Q�P���oA��Ŕɘ�ڋM[[��M�3Ǵ���?���z%�7f��+LTuk�z��dT͝�R�쐝�ͷ���s�e9coq��p⇶�	:������١_�Z|�ݍ֩S�/�����z���ĔSS`»9Z��#Q}�u"�z9gg^��|�����)V�ydⴝ���^���GYY�rC�Iʆ�n%�Ω,,�no]Ϸ�<�S+}^b�|	 z����}��1�2��;���M�e2�l���5$�R)"�� ��e����� ;�\<?�L��Hٲ�H!�V�#M���n����I2��/sss��M����:-�O>$�Ot����ft��iȌX�:����EHdFH��߫]m�ί�~�tKqk��2��������]P�@�ɟ)��i�>X����K@���i�3�+2�oEE�g��T�[ĤjV�зl�KP�AňŖ�w엖7X�XwMŤ�����7�*aٙ��}9�W Mn[�	�#w�_ʪ�Prr��i�_��&ԉ�z�$��(�A!.#���C�2/;�k^c��;I��
�xvɃO~�������ш'�dӹ�(��2o�7nZ�����-��lH[��g��6���
�ژE=Jw�| 2H������#��ϣ�}���ӡ���/�I7�q@J���! >o�h�ir�������Y�=���._(ę�7�J ����N��F�+l����p�nұ�͑�Dt�R
:��q��fw.6{�#��Ug��*���]�cY��N�!�pM6��v��۴���C,6{�0����)�B@I$c0��!�:9i�� #IǪ��H��5h� fkk���@ְo�}����TW���w{�	uqԘ�ǁq���O�jo��-7�*Q{�?�
d�_�9/� �y8����aݏѢ�Pq��'{ER/V&��xԶ;_H�O=�Kvѳ@�T�
���|��a��nVM�������$�CT2�י�N#egG�!<ݢ.űA_�/�U#��u�AO���Y���SE ��G�5�QǢ�d���;�FH�]7����԰����-Q��]i�<�������9�y��~����n��N%�T��0�DN���v�k�~���\'�O� �C6����T��$�G���u:#��Kk�ڿ`RJ1^�Y��ǣlF��TR���Y,6�����s8�rd������w��E����,�/�%����*A�jg����)�h��dy�v�g����"Ź �,6��֕������!��'�%��V�c8A;�S�.�A���踹���O6��懸����Y�t׾�F���[Nh��!/��y؊ͩh��3����h٭�����y��3����;�̬� �ߘ�?�/����S�5|��ʺhko�l0ML�0��a%����%����Ƈ1J6�$yb�*�t�. �w0
Ȋ-�i�HK�z�D�('R�Ϣ��a���<��T%�}��C����pu��b��X<<<�>~�pn��U�d*ܩw��G-���ʦ��FI身^u+�gYp���>J���G=�eaa���_�&�Tob@=���4un{�a��[X�Sۣ3����B*��^��@��VQV�s�T2}�|�ŉ!%�����v����T�8���0�a�S��P��5�)q(F��.�Kh{+��=`����(��R	���WM6b~�3>�����~����xC��E�uM_l~G3F�|�?��Kj��fo�@�����5�|��I��0q�*��S��Z˭8�ۏe�������G��
^#��[���f�D��Rh�N�@��o@�'[=zeF��S�����}K!?Xz�����`_��k}}=�*�n�f%M�9Dӛi���{nz���m�r� �%Y/X�$��s^���d��M��Q����[o��.��r��ϋ1�&��kh�����\�(�<=������ K�k|ŀ�G�c���5�Q�(�0�|)��"�	
��,��Iim�
*kɽ�Z�Ȁ5�dX>��S�-�A�[0U�8<��YU7	
y���WG��S�tv�l��z�/�R�8>�O���S^H��8xLt�Y9���g��3�ٶ%:�4)�`̮>YAt}�.�U�ɐ����]K���������AO�)ϝ0z�eFM���
:��������{�����|�g����c�f�z��W���n��x�Ju��^^I":�H�O�x��<YR��Q��^f�+qEV��~�� �榴�&bu���1�y`o�ly�ٔ�K�^��ωiOooai�Ў�R~��(3�:�O}�
��i�	��B��Duibh�$R�e��ڿ�eRj����\w��y(�}�%I�[Rbc�w�F��ۘ[XX������$cǞ��	*�8<RP���$�ÚޤJW.��%�N*�qh��+n�H�۟Q��^l/�}2���ETbӧ䇑����G���R�����m��11*�	�A(fqdF����������^y�s���y�*��T�Ј��a����6U����yC��H��]�aw(��ۆ�:;\T�7����<J�i�L��c�â|��D:����n����i	����S�����D��;�XX�w���w����>;�̉�>s���g*xq"��9�Ϲ��wY�ː�u�|��;�s{mS���]*)�X��6h���*�Xޟy=���+�UTw��mRet�3��12B��4���^6�/�(�GpJ�q��{X�b���|�Cp���&qu���b���7�2A�ʧ�n^����2L�:�����)���Za��訰Di��a�8>OMLH3�͔`�g���Xm"Q9�Tj��J�jj(����)
��401Z�+-��Pq%��,��A{x:j���ע�RL�sVz�
	'���e���$ҩ���[���(�5�]�j����ʣ����R&�Q?��</k���ʽ/5�Tg@��(���̮(7���0�d���0DgoQJ��6�$��?ʦ���Bh���>9�Qi)�]�pr�G�g����B�H�()�|�IUN1-jKfڡ5�c2R�w��}�����p�g[~��=Z՗��ߑ?�?��Hg ���ә�=d�Βfs��@u��j,�x�6�q�*)�+��V:�s�D^��a�ֻ�pwǽ�(�gl�P�	bh�8�>�&�@\w���&������d2]7��Z,[>�#�>a	���|��3�9m
<]=/u����+P	���`?��^�5-iꤝ����&3�l?C?���}���B�E�>�1�'�x � Ӷ��I�u�e�*�����i�5bIO܌��'�9�Y�%��I��iqG��"_�T�7�a�#��
�>�I}�oeDq���M��~4�s�	��¸v���'�����?�߰�g���l��P�����+���tL6���L���ȂT"�Q$ ޚk���S�r��v��ϳ��G�-z$�����[����C�?*�D둸{����(]�������(�F�-�"�6�_Ä_�l��I);,^:6#*�(�
�;�i@��FH�f	E�?pc�@91�}����E�N��W��JH��e��M��0�	I�Z��t�"��.�%}�j�a@��A��.��
�hT���1��N�/S���ٖ� ���n@G����>��������{%�	���V&�� |\6�GR�%>۳L���؃T@�8>⑨��8)^�i��:/��fń	"cK�J����w?l�JD�2u�޿3��R ����~C�.I�?�c��}����h���̻�dHY+Βt���9ww��3 ��e��tG(6��;?�H��Tq�����+����N���3��tޢ�l_mV�wO'kԏ��9��p��sS��< \��p�{�p�K|����G[5�ހ��7�fY�"����x�~3yF5�Z��.�ǰ�ŧl� �T�"���z�f/}��F#���fW\p�.�H@SE��U3��W�$��_�֞3���؇�{���L����WC�H����VY�6�d�*�r '�]g����5����3��_���G�` �b�M���;I�-����~�%��O�&�����O,T�q(⾏,="��Od\:��J󥦭V��".����Z�}�s�A�/A�s�+aE�A{=^e6eQ� �%.;��e?����Z���� J>���;m9x�@s29�-���������:O�]y8��x�+$��(�o�������7�ងܢi3�K
��i���ՎE���������.4�AɊ�n>�a�ܖq���!I�!�K��ZURVf�z�l�g �C+��J��x��)3&��ʬ���w���:�e�h
�c�� .d���9aa���(�"�(�^[��,��a
�m�ٓ�Z"(	P�=�ҳ=~�)F��]n���G�|��N"�f8�xς����2��~��b��G͛�J��Z�Z&�'(bx]�&�R"�Y����h�� ��sRuCOQLyב����m��#G�e��=�Ԝ{��֝�kT���)e�&�}n�|W�c�W�����<��Z@q�^�c�|B��̙��S���t����E�O*�����i���廕��#l�k�R8��x-��d�/����yv�Bh]S����#.n:{Kg��L���4Л��cDk2���Eb$�*�Ah��t������I`o�qu�����]4������>���2r]�׌������M�Z-�G��f^��#%�z1^�(V�;�S��Q�,3����;�vIbi��NEh?�ؓ��,��p���n7�ML�١�::�~��w x����z�pa�h����(���v��G��p�rÕ����犦��$*&�/�$%�$��-�x�[
EK�R�����\h]�5q���(/Z�9�ĬDu�	�;ГD����
�$m��<��(Hg��M,��*�t����b�{u4C�R��Y8k��'��֮�k������v����3t�ƞ#�&w�=����&���^mv
̴Ż;��\�Hi6� ,yr�C,�����隼?��v�k��W0t%�ʹ�>�ֶ�d�Yo�����3��?�9�{�ViFZ�h!�i@EG�7̽��й���]3&���]�!�S���/c����X��|�c���l�˛T �f��p��c(�z�|�L��A���Ƕ�M���sU����&*��2�?4_`�S�@�#��f���o�ilD�]u8���ժ���+;|��CO���$���N�-qNWJ:��ȴٸ�ub��S�9h ��t�_Q<��.F�|Z�\�70�'�x�g^e�G�g+A��_Wx���[����d+�h}�`.Txb>(��'y�by=l�4+<��9׾D�Pgt�8Vi�Dۑ���Vi�610[q���}�O�=�4�����P�t���!U�8GxA+��H�{IG��AuQe˵d�c���%����w~�������,p��sM���w��w�s�:�h3���E���Q�0"���xI9�Dv��IU��q�����s/� B#���`W�Jm��@�B��U5:zB��7b�'�4���y~9wW���_.��Q5M�����MO�~�ƭLL��d,�=�����oxӝrо09����	_�F�ՌUX�0�M%=�O� �|�R`�+@�&�G�N�k���*{�Ӄ����b��J4����I��kh���,��۽���!6�jLS�<�t%���?۵�c�>�G���>�����x�u�I�NՂ-��,�q����:�L�x�6G�oX��2�Vj�����ڐ?\���y#���=�n�p�U��!�hX8/��S)ԍ�B鲩b���I!�H��K�1�:�q�[QP:�a�\�����e_'=��+W�1�Q60P��F�������T9�01�`���N''�F2�YS��&����}�YE���X���}fU_�	1_�u�zߛ6=o�e:�9	>+�v�;r�Wq`�X�V\���b�{_����������"��Qƒ���fb��5�PWW����)��������7W��iI�{N���0�e"�E�UVi/ͯ:\���m��r��0�noo)��e�r�-D�G�s���O�U�a-{�AD�k��yL�ّz�'>5H@�M�1.�&0�g�
Z�ݝ[S����h<��h�<x��m;N.)��A���:����*�3h<������5a�tu���F��Y|��7j��nڭ�.�W�[��$P����Y���S;ׁ���ەfi�i�ɒ�����~[��yd�a�r.-4��l����ȑ@J�b�x�V�0����4��$][��ZÆC �S�d�\�[]�p���_ŭ�r�����m��ټ)�x_^.����9�����V���?W~Ć/h�՞��1��_�o-��|=H����8��8o6,T����қ�N����tW"�W��j�Y��i��>������<�ͣEh��{ي�|uq��#�7��������^��^ �����|�ep��XdL�{{Y�&�!�C!�7��r��������9� ��m{T⟳�1 �T!��l<Ȇ���O���
�6��\l8�V�wd뢒������k�Z������o��)u��6�e]�pJL�Z�C��DN���:����L9q��wR�n�!+� Ɋ��o{�kF�P���h�.�<�Z�ök���=���/�!�l��G�Q��	O�}�?��I��m���n����U+r�������>�",���g�I���`Vμ�������M��/0�8 �5���C~X�щ�	��	���Um�Κ�@z���Ӻ�B(h�%�|��>�+�����>��@�}�����j$�K읨iqa�k�D�0��2Sszs�o_7�P��z�
yM��E����'S�*7��L@��Zk����;�?�ny��~���f���o`Ň�H�^|��� ���P��*g��A��yy���o�	�gYV k��4�ip���m\3���d���W�)��0\�{ӜZ1�����*6;6���r�v�T��S9�g[CȎe	lD_،���G4�:ǩ�rM}K�>@���,r'�E�\�����X�)�˒z�;�~�����^D�4�T��+�-��3WE�;H)+�|@Bcg۷����\��h�r�-���K6��w�Xă:m/f��rs{�B�. ���5��Jy���D����&���I?�nk�C�{lR
�U8C��}UC� ���fU��y~+y���ZTSyT�A	,�qo~k�t�-�zi/i��3���%'ٰGU����d-�GUg���a=�M�H�H=X��_T�|�-5�q�k���}�c�ʅJ�|$o*�g5��K��9}��?֡Y��ӈ��gyV��86cu���=�q�����͕	;�� K<�>�Y�At{|�y��[��/NJ�B�����2��Ϫ;�]����! _n���Sp�j���s�'n,���u~�M]sܘt��>�t$^�C���;���zmC�\.���(b>C�.>^o�0��B��*6����)�H.qބ�r9�oM��W�N���#�w�X��T�Ywnu4�HO���0gB^�gU�/��4�bԣ�+�Y�0�������ztL���l<����+���g���0�%~s��k�|��c��]1����(0�`V�K��k�x�,G���N�9��������0ơ����Q�v��V���YL$c�� 97�㳍�b���o�'e�xWY�"�aa�|O��|�����fF��O)���b��"�7�Zw�2���B�D�oEz��q*'3N�p���	��6�T�8��ʩ.Ih��|���C�O�ǤsN�JC�a�"٤q�
G#�?ay�-^J���O�a���P��J\��:��,^Ϸٗ�̽�C�&P}����4-�v�_�@Q(d�ey�=)������I=o���3N�Kc2'�5�	�?g�G�&..���m\�Cռ�-7���4=��%n���UcN��������b�����%�I�����/]�e])z��qL1r{�r���d,U�Ȟ���~��v�u(q��$z�Ԝ�6c
����ܲ\�`�W���TY�+������� �T�މ���~���� ���J����}��xh"���8R˝���8���]�_/e��"EU�/�}?��S�&ǧ���M��;���>��B���8r)��8{Ɲb2���ݹ\i�����RHt7�Qs�����U�4�cFI@(5k��5�ħ�n�s�.Z.5��;U2h��<s��'(5­|�$J �㮝x��肎d�?�7����So������@E�>ݟ���ݳ)o�j�րl����hK�ֈ�vkkji�A��ܪ07>a++��+�f���O�vi���
�U��J�\�f_�w8���W���h��(p"�#��������֠>:*6Ԑ��%���	+0G���ٚŎ�cF��iQ���m}?^��u4xT��"ʆ�ZZn2$���B ż����+���7��յ1�1���mAg�2AZ��}��&'����K��:z4��ĥ��L���~��,�K�����[!��^�>Z�RS�G�l�������@�T����40���+abb�Q�!�϶���hT䞜��?2��"�@�����Y�W&G��u@�/�+�����������"ݯa��~��܀��6Ut�8��\��~�O���������q���*��7���a��>Q��"���q206X�x�\�@�1}Zu����NչqB�O�]��hԻ\�qd�0ݴ:���\|����e��=jSW/(,Y\�9�ifЊ+S�������N�Z^���E
1�|ju��r;�8�^-Umk�l�`�U���֞#��Vo���Q�꿾D<�6��2y��7���*�>%,0:��y�`���V�es^u�����	�O�f��g*�]�r���n|oe�O[n��~�R����	e/�x|i)bl/???P�:��j޶>Ny���GP2��<k\�BEu19�j��8IZ!=����
AY��m��� �>>c��v�0�� *\�fEaII��@��ܜ��q��J/]�A����u�_�z�ް���$e�<�rqǉG��S�Y��Ic��䕛��6D?xttd�_�a�=���U[5z网Jߓ�*,d��!T	jf�o�I��;�v�v+!�6ڧ�����P��D�[
}�g��$���ۮa+�����l]8-=]��*Ƒ���\��P�Cd�'"X�TSIE/�j��OM#�V�;���=^ܩ�^�ҿ~st��?͗�v ��}u�jf��c*��e���|��T7Kk\%�W��9)�|����S��P�"���7���ʬ��}��2�5�F�t�)��*z�\�t�߻}_�	h�	���,	����Lr��d��XVl��QV�^��]l������l�L�9�!��l�)����vC6:��h�ʷC����n�`�-Y�կ�D�<��DU�����w>b�_\�>��˛.�x��M��u�(h,)�z����f��k�f_���9�ѵi��!�87�:�����������k��"��ea��BKL�u�N;�/w�/Ld@|�f������'G�v@��{���n�!J���L\��u%��vd�����}�w�����^7�U�R ���{;rJR�PTKhoI��!��>��&=����m2� ��VU|&V���Ƨ���KII���"��N93�C����S2O�M�?P>���W��3����G���ܫaaaU�_���+'��O�l0H�r[�\�5�-��>�Αk�*��Hp�U�EAX�ЬF�L�2[�H��Ĵ���"F��s,�7�ew�{�t)L��1Z@��r aH�E�$8UGG��b�j��[��Jm�������s�H8�]_;N�Ƨ��r���'e�r���?�s��ζhYht$o��@��*�K	��yI)�L���O���(ZՕ~[,B�Cgs���Z���އ�{\k��K�sv��8�.-}/p�t)n;	���B1���
��������TV�8i�U�@�5c9�Sz;X10��9����S������p�U�c��5p#��Ob����F�9�g�n_�?���(�q��O����A`�7��EMN!j�n>2�YX��~��2���=x�r~�y�b�A��8eKs�^X�l�������oĨ��wEl8�NQ��'���Ͼ��%x�侣�{�C]4<����[�zBѶ�y~Q3�n�φ_�FG��B���-�/��^V{h�h�<	�U��Ȧ�`��d�t���HpE:'�&��*��x��qdx��y=�\"1SY:�i�c����^��>��ɭ+��U��bg��ZT����b` �] /+.������\��<iV�=R���eZn�=Lα��jؿ
yeQ������"L���Û������h�S��q��hמ�G� ]��\��qG��ToLC':B����Z����U2��5����T�08���|fZ��C�xEW���J�W�}��e�Ģy�K�w�˓�/�>%!1r�@����������k�yp���Q` �
	��OE�)[yP���Yd_�!�d!}��`��iV֞�9���R).K��<��k�0�w��"4c�@�O�=jj%3�_��9@�����"dM��}huab�t����M��ENif* �5����6}A:,�=�4�Y�&§cΜ��+����+�n����} c�S����
b�{�Gi6>�GA��K+ڋ�)��h����h��>Q�cLAy������1!�mȢdc֘��Fӵd�7�&+�`�	?U;�N�۽cM��g�E4���/�1>���<y�c����g�M����}�@I}�a�7�d ������ޯ��T!׎��jO��E����F�J-��� h}��37zSF���Qo-�;澗�|b��|0yKo�QRRbik��Uv'V�tj\�:�k	��O�a&	�$I�����C�5��jv�^Z�\�r���f�|�W����&�Π�b,�<��Ʈ��g�5e2WE�_|T-�@�čz��*�g��|��Y�bڤI2:���U��<�G��4V�YTy�wK15>3KPť���B�bj��¹���-�Y�Y�q�B��9�W�k���5��_('ݤR��|t��Quf�/��Z�u�.�-�q?c�?�k���{c���/G����;��C�JK��c�)�W��WQ'� �R�沛i?�<>�7/!���"�x�3�㾻�����l5bII��P�{��5--�K�n����J�}���Iq��f<@��D��᠊O9خFZ�m/���Q�'�}ji���5�Ս�����C�<'���?�c;�T]�2s��g�mT��Lu�g�ч�/jB�vv�r�9F,U:�pξ��g	w


�LNn-!�G�����W���,A$�~l��K�NØ���3dE�9D�1�5����*m�{<��ʆ�Q6YL��{��p���;5���B+S���q����c,���s�-�ZSii��l-v���������ܣ�H��MnCn���3ꤪ��o�ٯiR��2������C0pw���l�c*�5�4}� 	
���y����"����?4���:��DD�4r�W���z��)A���S��IU; �/���ԈVI٘�6];�|�Դ�ymu?VWW��*JK���9�阊l-Z�S<ɉ%�FyF�1"�6�"�^
�@��=�Hv�нe��~&�%���lX�6�	a��!�A�>��]���=�X�^$=n�9���n��]�؛��fE��=��v��ɜ5�S(b`+H$�^�Mp9��UY��V:hļ��deEd�%�E������s\~�w�z�;��U��EI�ֵ���[�,?`>Ҽ�4@H���-��GyMi�i�[��0�ϡ�՚**=6�4�s�����6�a8!P����Q=+!Ų�qO��֔�H�}�߉
A��R�����	`�T<��Ѯ��cMQ��M�1ɶf$�'F�Q�^�ԡ�<�=(JÇM).4@�A�z�g�89���ղ�9o=��z�24-++�����7gM�K��#���R�U�x���V{E��=K{A��5j�D�Μ�T)� %4_�Y��s��+:�d�<��)P�z���$��n"}1�u�MU�~����{�8[{�jOW�zrބCgȲ@9�\׀V<���#o�^��{YM�V?����7/њj|�5&a3�j���M�<a���y��m��;K>���3[���H]��<+�.��Ň�OW���,���2����X~oX�8_{:�B;eK��n%)<>Xp�;|C(�����%��� �g����l4��~��C#�����&��o�� �?��ͫ���=�� �5r���:��J�O�zQa�ȧ�Ω�F_]��1�_�[��fg�d�����2僒���j�6�")��EF�lʹ�\����	Q!�����M~7f��AuX��`�Bg��>��Q�K!��ri���q���������o#p(c�Q7a3�K���לWL~���y��R��Z�y�6���[�6���ۉK�@4�"�V4�p��|�#ܑh�|	�
���|��a��y}2�,�J��\X[��D��c4TD�Lc����ծe�B2'{�gҠxp3�q2�nb�2����y������br��N������$���@e dSK1w��R��z�G<�ֲ�������>ř��-�±���l�������Q��?=���<蠾r��B&
����;>36�����g��h��$��~|��.z5������ǡ���&��~�7����]�y���NS�֍-���^������IK�Z�&'��8�v�F��@-��swp߯�d�_����nk���i�O	�%�'���夭�l�̜K4����:����#UQ�#""b�~�n����^�S�1I����~�@K�����'s�"�W �T��&p�ۍK;m@�D�$��ǣ[z'=\C��E�{>�k�'����+�4����L�85���1ױ���);�9�g����	ݖ���^������w�R9����l��jee/�n�)e��ef��$V�[�a?^��S���ʨ3�^�es���-!�I�p�`l�u�c���K+a:�^�@�>��Λ��!d蛽�M�J��n5����B��M���j�n8�.�����4&F�\D�U�I8����V��뷖!��	�K���lg'���U��AQ��9&'�Y`�/+./W�v��
��`����ر޿��'*(���n�RSS�?�"&xXZ>���U5�Bz|g�Մ��~&�ov=u`<��KgD�^�7c-�q`�lb����z@��˰�ӌ��c�,�_. ���QYcEsxu���){�z`����]S�G^^ދ#����;e����� /M{|����n�`�}�K��]Q]���0�� ��s9�*9���/�j�T��3]W\TuJҟs�P2]��3f9�+C�cE��k$w^�a3��|�o����,!�%��^�G@u�W�d�n�}�ާNAY�Y7�T��� ��G��9��ob��._@J��a������㎡��Tk���{�טB�9�F�AZLZ�������YYY�jl��=buO���N�N+�X[S|Ǟ��bٺw &���>%Iz�ʎ�@��~{(ѣ�����y{Y�+Ư�$RApZ��_> e�f���c�p�	�X��[d�vI��=�"��~gd{�В��=S12n���="`��Ah�e�'��K�C�೓�5�����<l�!���ˍq/)Vj����9�%%Ş��񙙄$=q!Ƒo'KJh��k�}%�|V��Q������B���_
����,r�X�NOsS���,�阈�9�O>[?����y2�*dv?�b�ƐP9ށƛO�y�4��Ot�^�qlf��sА�Z­�=h�6�[>��N����&�>^�~�dG�l1�-ӕ��עǙ���gF�!T��w��9�߉��X�4�)���<٘p>}�Q�o�!�������捗@wO�b׌_�E�UL��s��k��e�������L����d�.IA�Ӫ��'`����J�Z�}�z�R:��^:�P֊f6�Tڮ�sY%:�K�'GqOz`����8��_�$���'����^��y���)M�=w���U�]h��ì��#)	g����MSIA,�i��K�@=�2vD}�lҿ˝(4%�-r��[��NUl' ߳�H��Ʌ��
�9ݿ^h�r/Jݺ������QBBb%�(+r=5[�j�����nP	��1~u5ώL�S�$�?<:x8�8h�r���|�E=���0��;B�Yʧ��K��33P���h�^���z�E���*��͸��1z��ȇ�ӕ�W���Vi�	�>/�7҄�U3���+��KJ�]]]!
zq��`���$n�C�fa����KB�hኂI�� �*�aı4D���+�eo�z�TulX�g���)��|J�|��ܻ��Ҏ��!*��M\�o���5��ᗸ�������偳��R	�2�J�K$��]Z����ܬ��.���H�9���q���cc+���%�
|{10�������G���N 5�3��;gv5��(�P�s�Ϙ`%U�`c����Nc��H�
ka�T��S����.];V1N�8��ޯ�0�ڀ� ���FSK�j�?�X�=�A�Uu��iU1�Iw��U����#�1�l����U{�x�Ӝ���v@�ĝ�u�@��z��\�	%���=���W�=�϶�U�0�TR�c���8�X�~�� !��f/w^��г�f����ե�ⴤWc�Ny5�h^�U��#�:�]��j���ŵ0��΄�ڔD���?ˮ�k<�UޥiI�p��q�����lޔ�g�yޔ������s�ٯ���9a!Hְ[GU"�q׍n��_I��&��%���,=x�q@�	!�kиۄ8d#����U]��%�@�˻�Y}�n��]��?��#b|朮K#}�$�m˩)�I�H��m�t��i����ւ6)ɴf���6�n�]����S�X@�dL��� �AܵVh>��5�-�
�A1�H�/��T2:�%3�4bkq����97�A*���L �Q��j�S ֚hJ�qbY.��[6x���>�¤����"�K�՝ތ���:����f�
���r}Y]]�����#n��r��Td����S�#�s2C�gt�����e�� 3����R�(�;���+��  =u�y�U��׬۪� c���N�Y4P'��]��s겮�KKd�g��>vfy�$RN�2|8���mh�}�!��I��9*�h���5t����-�����[�B��ؙZ�*JTq]���$�3V��Y�'��pp��m��"t��ͣX:5a�qW~���S��컊|J���3Z��F�����̦��m#z]��{"G�E5P�g��	T�ѵ,ð�����j��ˉ��_˱�Z#&��{�,�&���;�����l���y���<}���X���tS(1��S�M>�G���|i+H.m������CCK�V��������rܬs����
��,qx��IP���m��[VF�LB���fP!�1$$$� .W)�g@aS�>�fq'J�s�V'��֠�d�rlBi�����s?2���?�
�}˴�f�n�����6��[]ݭ��8�!RCQ���ҘE���a`.��#ź�k��L��oU3��^�\H���kR����_k�i��S��ϻ���KRUJ��6�ٔN���4&�}ӝ���p�~cf�wpv��j��łi���A|��m&;�HF�����IQt���mi��a�ܭ�d^C/4��\貞�kO���R� 1��x9s�MnH~K� �$q.�Z9ڭȜ�4LqF3)�n��Z�V�9B�_R,o��X��YC<��wh8ɓ��5���G9�|�ߚ����♶�r�˜���&.De�JK#���M���󌪴*l��Y��E9��Y�)�����U��Qd���ܱ"��`#>ף�*c�2u�3=!�
�V̉���	d�\�򢍝�`��:5Q3�v{�E;?��<���}�g޿t��G �Y�V4���<�X�!x���Xh77�K��F��9�cgo�v��������	*�]��T�b�h>B�_����z��iVi%
:u�dOےb���^Hf��'��xK�jW&��54�pL�g"L��>�.8g��{�흽^=��]Ǩ�(��O�P3������эfJ����I&ػH&ht��Q�iʍWx�vƑ��K2��#B�CU�^ rpp@�^L��Q�Q��O͌�k*��s����Ws��0��*��`S�������-_<Ӿ�ӧ�/frsD��g"z�������,d�2��0��B�cu�q�n#�_~��Ys�H�Q�z\�'��U�`C����j5e;]�7D!�*�8�"��GGe�k��x�������|u咘d�I�K�!���L��m"Z�m���E�l�;�Ϳ��<=���5c="�����:::R�JZ�_�� +bG� ��P���..��J"vuU�ϟ\�Εg��:�2��(R�	H���ߡ�/�*ӊ���=��O2�՝ ���O�ffW�5*��+=�h�J?�
�B�{��z��%�>Q$\ep'��2 �]zekC_f ��^/���dc���I�����F�R�m�����=a货�i����버}�\%��$<�O��
u:Q��|�.'{�lȁX��&r��Z�p��lJ�R�G)$E>�+�O��Z
����yN(y�5$|�[XЖ������|[PPP�S&%#s������kmm=>>՞�������ԓ��髊X�$LY����_�������		������QW����,��Pz��@�I~l�+LZ�h{I��n��I��d!,�90'���+�QH�
��w&�{:���8�ƺ���M'���%EE�	Q�..��_�U�X?��}v�� ­��\��*���*kl���������,.+����BX�� �Z�ik,D�9��EG~�qy�~���C
/���1���WF&G&j�����B#�X%LIE��%2�Ѫ��k��l�e��F���@�u)L$l�~�����-�����Y���(+e��go#ZY���ѤJA���AU1 �1%S'�V�H8@*���9��幦	�/�'�?��@*�_�de��h�Ø]��VP���ىN��y���2j�	�?�{����D��Ǐ8��}cP��e燥��kT3�M��/
~�hd������NN)_.;�`gyk�RL3s����KKb�|�b,���.�2�����5ؙ}�t��mɣM!���>���5�<�|�'���h�Z=�@�����H�\�ޑ332s��h�c��f�ܑc���d|��d3��?�	VZG_�ג�����s65�śC�h9h�b���7zvQV���#/mF��N ���eu�#a�%Wt��Q��楥�u�gF�VwB�UD�)P!w�Ө2��o�Y�+L�*�z�x�<zk�!TE��q~�
ك��|��m�F`f����ee�")|�m�h��+�\YɳH�jq\,?�[gh�{R��\dI���wne���А���U�R��.�"�a4~��$��s�g��i��|�,�;H����� ���̸�6d��}�p����Gj�m#HR����%���n���ް'p�04tKm��A�6d52��A�<�ilT�_������CP�[���ͱ3��pU%� �da+f�v�Q�C��Z��=e۸Nfz�E�b��J��Sʓ��.����ǈ��oP!��Ň�x�(���0��]iI��H>�0ԲqZT|�B�p���}_%!�5fms$������!��hkkk2C9�dZZ[�  ��?������3�
F	[�7}22c[! ���*I	}'Q�y��m������e"r"⹡�;?��@+?��P��/+�/G�ս3�쉵�	Q}F��Hǭ~eA"���y�B`Xr��a\�N�����7�~P�PF��֔0�BF���$�I�B�ƅ~M�L[տ>8y�N��I�xl/�g�o�,�H#(�Txg�K	Jn����-3An�����e T���� 4�0�!�@q
�@�2^ț�o�Z�\
I���V���bG
�� gZӟ�n^]x��Ў�y1�{S��-B�lY�Lat��D};!@J�]�É�@��Wo#�p�b]���B�P�	J :��;�l:�l
 ,���w��Wi��˟�� ��_ D�S���'���W)#�����V�U�!3����dx�TjAA��R :�gf��ofQi�_A������MKK�q��?c<c���WD"��jw}�4իC�W/�k+8���`�c8T���Al����B�8��jߙǁ0SC>{�5_6��-'(�����G��;�����a�Q�wi3�X��"f��=�����,u޺n��C�mд53��Qp�֛=p�SKnYi��F,�׉�"P/.�Ɔ���X�D�B��Nub7���T��f����G�i�F :�� ���k��|�2�I��S�B
����B�؜��x���̾��붖����vy�"o*f@q�D[�CgF�tA����~pW
��<6����yppP�˫u��X�3|�J4��4���87�&���-F���YM��,S�1Q�,67W\�O�i(y���Ș�H�CD��gi��	ކ+��+U���h:�$*P�}$�Z�ۑ�jd�9�H��L�L#/3X�IZT�K�P�ڤ��/_��ⱨB�G+ֿ5A��{$� |	r�%�����E
µ���LMpy�L30H-���_�_��!\@��>.7�5c��h�:w��~��hj�:U�XH�Э����g9�}�K�z92�WT<cݤ&#��vuu%%%�s95����3<�m��g0S�}^+�\74�.�ՓӖ�5��eG�4���'���K�Zt'u��bRB ����b��hPde��U��h�� ypp���	�o,��UUUߊD�o?���i?Ga��F�J���L�qk�Ƥ�4�Wk��'������jM˸ꂻ���6����'��� �vK!�e�]�Y/����-�ZII@�'�wQ�x�,cyQD(H�q�;wt��-ˊ���P]��������1�ʃm���Qc��$� �t&C�Ǿ"d�us9^ڳ^�8�6����y(���K��yH�A`�H���zֶY�*�{M�w
�WX*���w�$q�!߱���2<�Ikwv%����10��⚬0�]O��t0�v�E��^7	�N�Ew�5�-]�jߊ���(7�������2,���zqww���]B�,w'�;�-�܂�������w�|/��c���鮮:uNO���<�a�8Ggq�'��|v܇�g8X�E���H��ޢ�K�����h�E��N�G�?������y1�9���g'4���_�Z"�����k�������*P�R� �.o����y�ĩ5�̑�u���T>��d�E��5w� z�2V��_8����V޼��_~��f�{�����̔7fC�+;�m'����{3��Ks�8\�J+wk�Ǜ�r�M������?XB4*��բ^���hWp��Y+��� |��\����7�1���z q�8<��kSm�Z�߃�0O�Y�OD�Yg�Sl:��u��(�p�K.>�A�95�P濭�A��<�fd��b�J�j��ʚ���!yF����k�P��;��\�W�1]v���S���T�G?B����&1���x��ѷ�����t#`zB忽��o�8�������rr_
0�Y�}���%@��q��<?T�ٞH��I/���R �o���m�K_w����hoAz^-U2���Lc"���ۤ�W�4�iR�\�~�����V���l��pzs���GE���n�%��vD�phR�6J�$��A�L%�|�7��'��xg�h�X��׬J�әaF���q�o�;��1a��p��i������e����s1,k	�����e�q�4�0�R��,[��)���hQSSw�VwZ�vY�t�s]ߙ�y	/��p�����	;;;kߨ�1Ο=�{���s��̽e$C5g�+�2W�op�Z��n �#��\�����?�AP��M�;�,V 7��;t�\��UR�����a�z��j̾;1*p9@��65���.�ů��)$(W&���f��)��W�,�����赳�#�9����d�d6������ٙ���-�n|�:�ɐ׻���0,aGZC#�[�'�9���{�[��"��<�J�HF��J�Y $)�k����יt`��'���%��;�c�B���)iia���e߿��~�y�%�!�K
t]��J`ǯ��̆=�,� �~"�5�����3:��y�yPx��%�����**JP���+��AW�3��'�9��|��������5w����r�v;���E�9�Q��n79G�]�I�Ɔ�=�9oW)��~ǲ�i�Sz0$k����}c���6��e����f Y\R�Ճ���cX�a�*"�<�z^�[� �s�%L�+%��4�"d7#666����W5X��H�s�D%���2��Թ;�鷔���}�� ��bC��㰾���E}�vڮe�+��J�Aۋ�����j���Qm��6,,>�������(R�ʀ��y���;������#�?/��S</����n![�z����Kf[y��A̕f�rX�F�����e������1�yN��p�k�e����r�]!��G��T	b�j�� �`���U��^:���`8�tjz���D[1T���Pŵ�*�s2S�^��"�@���~S|$��7�~EKUӶ��'/?_N@�C_�_|4;�_��)Ú���l�4$T��8V ��+o[G.GY�t�Q�ŭj��d6�fC�-|!��ߑZ�A�}o8���h�u��9!�^[KIN�Zq23�_�L��TІ��ڞ�_�!������ꍏ�KO� $����ی�c�R�Z�)�GZ����>��!j�Hȁ1?��j�Z�f7�ȅ�<KDoj��J���oM��o}5�s%:g���U�*8�������B���@-����Xr�8�Z��бX�����d��^����\�h֋=��
�����@���\[Ƙ����-\A��E���9��>�}`჈Y�q'�Kh�������n��X[3%���K2�z_\T��=\H0L�d�d�����d��aҬᆱ(֘�u[��cz�L��QYW�²!�d߽��������zx��p����.�zU�}h |!�4?�Uꆧ5�{����I����Z��=}����(_t�VoD�jQ��9=��)}~��!��zI0�z\����,�߻
$?�X��.l�'�3i�����~bZ\\��1�m��
q7��^^�~��.X*voĆ����IUL�½>]e�8�?*�X�'� u��K��a���J؟Ov�l]�нNQ!pW�tA�U�+���13	˛������4u��MGť�������i�b]��>��H��a�,#��t[2E(>>��*zz��:���5� �5:S4�P������y����ܭ�K�l��Ot[��������b�|8�aUvv��e���� �������|�0����Q���|���##�B�j�!q�u��]k�c�b"ߋ�����t���"�,3�j���H-*㹬�j��8��������xJ���9�@��V\�L'�,���.ohhi�L��H5��b���e���$�R��.���1[��j!9v����Н��m��%�
��"<.��ذ��=I��X�eS8L��O����CM��4�h��-'w�s�3��$V�/uZ�/0�y)����T���b���Qp�w�����#�TU��!g�pׁ���8����O�ICi����&�������W�\��lN=���G���a;�n�/X�e�55\*F�S@֚�� �T�1��Y0�R�< ��3ç-��H�v�0�gP��a_Ue�[E�m����pІ~^�URRR��.���sF�w�����j]4��Z�NJ�ҒA)S��R�ՐrDϗ�r�\��r���QlU���f,��bc�_��Q�p#
�\P��I+E�,��#�z�k�|wMNH���FGs=��/��4���1������F)�	�$�)�BUUUI�	(X(H���l2���%���1\�����U1�(UW���ǩ[(�I �̐��/!�c�ǈ`��G�P�4�`��%/u���bd�E f��?"<�Y���t�u����>L�b8Y�(o3y�N�<�l�,*�I@Y�
�y��<tq�Xmf˖*��TE�J&���R��BB�Nq�o�U��%���E��<�Q@}�i�R �_Oe%Qj͉C��t4��U���������Z �"����[2{|X����/4Ur���^�Ar�Y<���YKN
0T.X��*U��/���Q̹A��c9x�� ��
/v��1ji�B;�X>f���ٽP�/�rzS ���p�j�&�3ʳZ�Z���_ɞ�`?��G�,���CIfH���E�j�Gr�p]�^k9����zu�a��闧�����ot��O��(��ln׋f9g��>`y-�K�O>�l��#ϲ�:貒vU�m�I�>���nq��޾�H�TRٮ"�)�����D ����w-6��m��?(�		)3���3Q���|�r��$�>_�u�)�n����Ct�������"�ᗪ3�X:��=x	ӯ؞kt"λ�$+̸}������y�(�eG���	LӪ-�$��%ǁ٭.׶�����3�5/�;l��/�X��p�7�2h�==T2M>"K�N|䁱1i9@�]Ʀ�л"�H'6�������=.qI��0\�� ?@��Q5{{�*�r������� )+ii�hAܜHXV~~���VR4�zAq�䖖�BƉ���]%��B�rA�>Y�^0�e�~���,͸l5����.͟/󉗖���N��7��I���Ze�B-����LDt��
�(+����|B�U}`8_�H��h;��sY�
~���äE��qvfF=H�!R�G�S ����L�d��Z�:�!@�k�@���Х��&�A��CC�US����襅~g+���2�[����0JK�*4O���`5�	��������6�����A�\�c�����T��Y�}t����K	����U��I ��"���F�5O)o|O�WT�~HC��2ܜ���)����d�E2�gL!���櫓��Fo�K�5��~��8��ସ�Ӓ���%��OB�r0�Q`���x+��$��3(N�������@�J7�S/�O�MG����hCfd���^���5����tuU�{.��ɔoN���IIIᤜ�VV����m�V��2��{�XtЅL�Vm_>Q¾���frR����#�X� 	%Ę��Zo�@��P$򫈌U�r�)��ht~�jюRN����RZS��1j�ϟҗ�)����#<:hNA���SS�ظ�⹓���,�ƿ��0ab-`9ń��ͽ�ۇ �cgq�ݞK�rR��_�h0��j~^�Z��Ii�c�n�2}���Bu���ō(�?(���|x��'9<��5���u'ѻG@��{���L2N��B���m*������A9r��k�q�@�J�w�5i�I>��T��$��N���G�qq���@B:L��}Ʒ�ByR��u�.�cr�����p�yo�_�	�縇�S1�Y������ѧ��=U���e���,$�n�C��i����T
��Ta�+C������T�Ey#�P)�9^K4W�/�f.���tg�"|Br�矝ʤ��_���A�k��0�{~᮶�olmo�{`�Q����s�s 9��hSȇ�e�Y��aB11x�?����CH'l�2��Z�^�ѭ ��Cz�/SɌ^H@	)��w;޲AJ,v�6hC�������A�#�Q	uf�U�v,C�>�IB��4ͪ"������_�����Wyr�&�������BI��R�v/ܤ������*����S����ٟ|D ��]LkЪ[A�U������������w������  \���%m�B,�#%�T'��7�;��h"�{�$%�W�-��2-W�������������~_O/fd\�u=�r�a'S�) &��� 8q'��.��Ƨ�-S��^8��|LhT���A
���ϩi�3��R>�B�g�K?�,5�m���{^�
g�٪`�"B�yU���t>j�-�Y��?,�+)��NV:ꀟ�� �����(���~J���SyE6���<{9ި���Ω�J9ko__�cm��;~��ɄK���:`g)>�%��el���F���R�YqM�Yg+�SOK����:�A��5圾FǦ���0���OII\���M�Ū ��e����&x�<�qJa��L
������wᨕ��fcA�t"��b�{埽�u�m�]���!L�<�.��H����B�ES� ��aW���ؽ�go+B�z�����5>]	{l�{�&S����kx,fx�\y�Ϧ�.0�y���u6G��t�:�ek�qp��\$�*i�퀀��8e(���ziiI2�1�J&Z�Bpd:�;t���5[l�2���e���K�?�\k����:Plr���]�W3/��ME;�ڡ���3k�(h)�3ghP��/b�tw��P^J��Y�Y#h�y��֊�������3�>����'�	Ow�	R@TԄb*�h�F�"�@xqr����)�պ0���^���A&&*�#�y�7�;�[��jz
�Yi�����ׂ�\�:G��`�鋯ɰ�SW04�ٽ!e	견�}��v���m<G��;?Ԝ����9R\�ڐ]B��'��X��q7Z�׺���v���<��i�cUp����CÁ��Z+�GejZq^;���5ē�T�LN��ܙ:%����t2��w.4����"�9��{���Hg����@R�[�.�LSk�d}����q��7%�}]�_h8D^�m�y��88��<o���vh���QM43m:�[�g�Us�n���n)��;s�n5�{�c���Џ�������w��ɧ�P�xR���:�s��T��V��� ��y|K.y+�7���r�:ؤhDQ��_�� z2���,�%���+�Xq�~��>�WW�ۋIe���C��_^R���Ǥ��@��q_i�e�F�����C���
���Q�D|�Ֆ�������Ջv��/Yw�W��x/�O�����a��R���(p���z���������� _y��k��^�a�"h�K��x��2Y�;��&&�zڈg�ӁCD ��}�l�wR�u�&
I��u��h ��
@��y $����:j�ȼkZ�~LL�jC�C��{����_XUut=�V븟&���}��K���FY���d�2~>f������Cܟ�����ك��(^���u{���T��īp�6b���q�����&��&*5w�sR��?�%�գ�}�O�19����8��,$�R�=zL�f�ɒ�f�g�Q f��쳭/��W��w,���.-��3�5@ٜ��;��Py�MSگ�*c�[9���Γ�~Xov�⽩	����c�����"�pxh�{�0Wzx�#++z?W6���#�c5wI@w����l���y�^W��4��GK��)������㬬'qTuιG���.b��WI�	��_�0���y}�|3n���q��˽uPvE��mJ�J�(�_k�d4L��I��js��ݗ���?����̽:lh9l�iw

*WP�M�b��3"`��UZشT�͵fW�WG�=��x�҂Y��O[����X�q��t��A\ k�"�DFLG	�Q�g�h6�7W�:~�B����������9�"RSdϠiWѻNx'�F��E(�1tY�Ym9#�>D1���Ml������O�n֠&t���F�&��XaM�	�|�A���BB� tH5�}�	VM��)��\���䆰z�nc�_��<'χ�����΄A'67��p��8���k̟�9UV@b8k�r��ac҂ȅ�Z=3b���v�MyJ��N�i�#�E/++l�'��� ��|�9�A 'A��x}n� �&�߶����2J�m'I+���kY�ʃ; E���+��is���<[�.�5�]�������8�A:��

Rv+�!ii�;{{C��=.;����fgs��a����	�us��� �)=
�{�4Ԡ���B��I�<��Kpx��]. ������n
�� ��"�:ba�{w�LF�*�[�r�HIGGN�c���[շ�I�2���>L_�YB`T����0~���PM��خ}u������_�
��b�<�ƉfS���opU�'[��ݓ���epI9��U+��)n���PCl9;^Y�Q?�i$ŵ�GpM�E�O93���k��E�׋�O���s����gk؊��QB�V��w�F�����n7��������Z5�uu����|oc6v�ә/ٟml�,Z��"jBbg��^V�!+�.�WO=�����V�V�7@�ݲ�4���xl0ma(�/���D�N���Ѻ����*$��]N��b����l�=�Z��sDɇ���b!v~�	��r��_g���O�h���'��2]�_�˝���}�Q03m4TU!�U���{}��a��K�I�<�oGl���7�J�R�(���Iq11艅�m�X\O����~H!5����������o�I�}Ƃ�i����{��pr��=��H��]O��*��"&.�"@ϵ�+��f�u���/뭾"�q�5���Ks���n��e4�'|V��	e���%{h����ȳ%��uB�L��'�Ͳ�[��Ȉ��{��C>i�S	��b�K��әU���0̔�x���݋�uʸFa#A�OZ���V�#/�Ŕ�g�������6(�H���ߥ�qJ�ʝ.T���
���u�u�F����!��'��Tnև�F�]���O�[?�mz1������Pe=.���j(G���":�dW�pP8Me��n����l��h���G@s��&=o�xK)3����s٭�����P���Vn��K7w�_9a�e2����03����)�������F�^vqq�[��*����`~w���n� v�����d��Pm�f�߹ � ͢�d��n�P04,�e�ù�T�2�QXd�����|����}�9��iݧy�j��q;�}����``[zH9��h�jq��'&	�|����$�V�y��0��ʃʺ�@w}S�W|�@EU'27�)]�����ع�͑4n� ��4��+���Ľ����ν��*�CU����^�w���̉��b������w ?k|��P0�e2
{:���\i1Mˤۂ_������$�U�����o��X��B��������1G����Ƃך��_�F�+꟎o��%l�R�A8���p=�v8]A 0��I���L��&|vk^ĄC�W��k�����&���>"6���)�G�F���t�ie�g$�<��yr�8�N8�Lc9���e��GDt=��2b����Yt��X�l^�dm��rģ~~HF�(*�IUL���J�y/,�a�������/���km�t歒�L%:���{Z�t�{�K*�H�j�u\����p�}y�=���H��V��x�]��	~5e�{��P	o����g�	ɿ�.
��("_"ኞ{x2w���l�*T&�5�k�{l
ۃ��֫�oYE��?n <���\
��(���@�}ǢI��$	f-��5�4�{�{t�b���V��� xVs&���x�=�Fj*��ce��*Q�N�.܃b����|��z3����å�����č��e���y�X�E.�������:��O��"ڕ
�B�����{|����T���݉]����S]m�Qz(�!�#".v����6���ʨ��K!W��a�/��kv�X���_���\O�MǿG��Q�������f��?ޏ�넛���B������]w��sV0tɴ3�1V���6�,/�i��@8�W��}刾F)m�[N�6D��O�r@0 ���@�M?��j����9Ϫ��,�qu���\�`�ʓ���K]]��-p_vSl��"R��v�2cN�Z�� T�i%�yvȊ���p=������fe�i��KC��={~� K�G��9e�)s���3'�f���j��Q�AEe��Y��v
�4�D+5 ����m#+��0��'�]�_Mb�7�kD��#����W�i��41�Y�}�V��qDQcH�ޞ������OstO@X0h��z��k����17�!�������g��U>�G�5�}b!.�^~��V����o�J�ìP �����Ϗ�y9�1}o�11�	<��K��x�C�`E���?�K���C���ͷ]��Z�^�L�
�����Q)S�8���:���x�B^�h��<�x��j&]��y�b����C�m�W$�͛�,�����O��0�f0�G��}:�q�14�7�K�i{�����M�t��U��쩰��]�v��H �t����]J*[�T<���zB0|'�=4*�5�fW��Ky����/��;��y H��>��U��ľ�9~�0Bܷ��u�HW�H��|.��<�~�21]�_�05С����{����hT���d�^.�TQ�`I@j�̲�-��3aA -���-������������S��mae%����G��q.�VP�8B�Sdsw5��?�9b�Dp��sb�9� �����#u|�&���_B��_�h�D n�A���õc?�;�?Q������v�����o�l0��\-W�J�������gAWq^O�y]#v����sG��W�Ec��,_�ӧ�NAb}X��F��|��[�UW�������筈r�I��=�G��6H�p��g���[�������;4_��x]ֆ[7�J�{��Q�-/u��-�] �B��.���ww)��(�E+��f>�M�f�  ���ҧ�����sbAXTv�5�љ"{�k�Z���;�_ק�.sL��s�ܲA $��Z�y=��&��-o{��bbWQ_���QD�%��/��3/�f��7�2]�OD3�hs����̼�&�F@���d��_�z@�� +.�����@:��_stJ�=j����w_�a�C��EPZʔ���lq�Ɇ/��3	�2@]�u?��י ��y��V"�f��ڬg��˶���}V��tA�/���m,,��E�(i�`q� ��(9(y8xnN�������)��-��p*1�q/=���'��/H@8��_�Ի���`�!� �B��x���*A���9ݧj��S
���o��ɼЫЄ�]�I8��c럇�$_�v��>=6
k2��h�灚/�`C,��3�/$K��q�{C��W�Ǯ�s��[����D��{/�����[g>p�C�l�:��On�z��R�7=X�#����3���m���v���(�6@]"�Q�z�5E��)_�ى%�#uO�{��	�Do�J�u?b.�Um�4[�d����M+�)��ɿ�m�߸��h��׮�yd}�x�d����zK�=�?p�f�����|��^�\�8�
�S�K�y�Kn�tHP�.뱋���O�++����~�ps�bT���":�b���Tl�p���Y(_��			)|K�O��781a;��=C�Y��Ut�\��o,�"����H�Q$��W�:�2we���N�=n|tz֯�øA���'�⤿���uX^f�.'�'�����%$�SWf�R� �7�T�an:[�g^.�=τR��@�5�4��J�����5�^bA����� ?�\�ٷ�I��S���x�޵{�U?�����Ѝh�9�Zj���tq1ziq����5���iէu�j+�tD��]�0k��4m�Y;�6s��a��䡇�7��H^N�u�z�CDiW�Ę�olc3	�neSc��xH����O�@8k�� LII�Z��]E���V��X���>��-��&�OD�/�@޾u���(4�����n/�[t��g�X�����4�!V;���7`�=��(G���1�k[�ǜ|�vg�_r(������Y9�޷��D%�Γ3?��AeIFbIf�m�	@�e?���m���R������0˚w=�]���ާ���a4S��_��8�_���o{Y�Ic��K��.�3�~t%�i�d
�}�e�$���}܎%-O��'y�/�y-���-�d��������ź��[�ت�Oe�Y��R��P�0��yyh/��X$��[�J�҇,�>A�:�Q�u5�vQ��?N�7�fx;F*
��܊�Z���%RSg�h �������5�u&�k��� *z��#i��a2�Q?Ha�y���J�pwR��2�I��u�0 9�����	��l��_���I@~I�Gڈª�S�	c)�L������GI״�?�R�K$�"L��m ��ճ{�J�`�����<��8�#���V�M�5�Y'���^?��^��[R*9��p^f,�{e�_Q.}��N�S�i�)������,���~���S.Y��y]����՛��1IzR��1�Kt
�5
/P��` ��|c�����1�Z�*e�a��T�6�'�m^���h4°�c(.��L\^��}���{ �x'�QD�%I.^v��5��:��`�8M����h�����	�clo��VO���\��wߝ�&~"b�buN�Qx�$��72�n�#6ow�A�O8�"]�����m0�Vj3DE��C��e].��I�F����j5�[�P:����r�f��sZ?T7ʏ�K*F($@*T�*��'�~����:�>�����`���+�.�g�9���jC���u���\�Sb�]n�o{�<�Q��2�նI�Ê>j��k�l�	f�~��5���H+u�HN��Ԧ�nB�bZPv'y/���ec�xito���}�W��P�1햄�EDD�@TgW�G��39���e�6�K-�Ou��5`�=\�_5�����#����FIAl&���\��^�Zq��蚸��?w����#�	�*��e��˔#��pex���=`d��߁���_�h�#&0�L��bo<ַ�h��z�»� @���Q��E�}���JR\@Z�_ "J�/���&+��bU�K)�t�@���/���Tϋ��J��ﵪ��LG�B�D �ڐ>*DX�K�������
���kEo~}�{��<�q&D���X����N:����H� &FW�֒s!(���8w�N�D5V���4
�G��F#���@PN�f�si"3iX�m"sf�X�D�7�Y\��l\*��VA���g=%���x�
�]v<ÙJ�{�fqϓ23���+��LL
J�߮�Pq�N����'�_��yQQ�v�J��O��w�K��;	�E}���-\�����;��NPx�������u�����:<��gFR��#^��Ug$DDR����U��3�H��f�p�c<�f��Di�0it糧K��S�0ăƔ繸)6�Y���k��1�ԉ��YUe�f�l �Cƺ��&��]V\��n6Ny}T�k���4-��u���oeLi���hx����U=�5t�����%������N�C����ߍ]:U/�rzbb��-,��j�arrW(�K �������j����B̝�1d*�,*���Ӳea�%wRRÉK��_`|u@u�\�݁1��驑�y�լ�k�l�(-�E�o�u�U;�C�`�����[t���w���.6%?��f�t׊Y]+ߊx0�a|�m�t?bEKnrRJ�����PK   bi�X�ة� � /   images/ca60ea1b-712d-4ba5-bcf0-f1dd45701dbf.png4Zct]]�Mnl'76۶��F�ƶm�qc�qc�N�_�o���>?�^{,̵�<gG*+J!������!�H��~�a``���_OF �̯�EUJ�f���LF\D����/�������zje ��} �,"
^K�v6:
6�q3:* �6�@|P��FED8a�K�AM鵷y
6�9�k�q˓��s4.�����{b�7�sR�������r�xm����	5���x=�$	VI��\Ҳ��L��6E����ZܘTIy�c��4n����bO�������'z�<�Q�w�ڹ�[�@��p���UܧJd��ʑ�T&���Ϝ�F�\�|��Q�Ώ�o��������M���NIg~�5-K�??�-����;��C�Y ʥ�W�8����xڋ��G�K)��Sq�U:	RBt�O���eP.��rΧ��3��nN�~�]�%���L����9g9~�@�a��z�Z,�'���[��"@�aW(5!��X���d����z�-3�c6�,��T������P+�);�0Bg��|a1�_`�@~���b����'�D<M��V 9����-��\��:�	Јh
Y�P�}��d��ƭ�;n�+[�Y�{��9�y8���Z�������^��lG�k�I���o�]W[N!p�]/�Ur>���I���,	� ��9v��/�^;)F� 1���u3�UT�_���#����������ڟ\��ܫ�8����͑�v�����{Mw�	�ם�㳹�qu�c�)`e��/6:Q���/zɮ���� L�p�<���,ב��v���G���ڹ!��G�'q����Z%Y��1�]��ޕ�r?�)��t-&��]�5���� r@��h�y)v�;�?r`�D46��U?�F��?"��hʧɲ�gl����bŲ������O� _� �ƣ�n�1�5��T�<���u����d�Bm��JGq5tj��Xl>�}3s ���ےB��<5O�e���HS�y?�>�-nw�n�2�S��~R�q���k��k�$	UT���n|�{;��5;�y��Ñg�
����,r�vc�ߠ�Cvχ��1�����ٸ=@Iĝ��Pb�.&a	ݫ�&���|��|�����6���P ��i����u04R��pM;��.*d"�T���b[�4Be�\`�G>���z��̓�����y~�:�h�Ϋ̅*�-��􄒈�S�u�Ɛ Ih[T�U%�w�+�'{~5p�?|��wv��Y��*�y�8���5�p�j�k��&x�i1�I'!"�C#��Q+M}�/�
Լ��js����a#3�]�+*i�4c%���
dLɱ�ط���[��Ϲ�QQ�z	��+w?�w�xyt-�if��ǆ�	�&CM2�Y�D�Z@�:�k+Z�F`�=�Y��Ώ��]�,�ޘj:,T.DVy���7���!AE=��u�D�&;���A������c����H�6L�T����f������}&�5:|��5��FF.����7z"c#�Q�vvfQ�}����W�g�"��q+�ϲ���[c������$.#��x��ސ���S6�jA�Qx	�@�rG"��R��{���S�U���x`���x���[�R��N�Qw�\�5Z�L�h>4
���/�%�x�7V�u� �,˝SFe���Å��� ���v���!|�-.�oE���?9]Պse� �\��찾�db�`̢|�M�A$�s�?O�	�gw���%�y��u�ʵ�s�ړ�1G/�f��?�q߮�#�OР����2�حg3V�!��`ȳ����tr*I+Hǰ��s�M��̮K�;8;f��:��u?��j^�q�F���'N-".���Z�o�`]|���s�Ƀ�F҄a�I�67��6d*�0
���r���5zT1�c&��~�B!O����L�`9h�SV�9'�T�<~��R��TEEERο)%ï�,
�������j�����j6���z�-lgK"�ڢ�"��n0��MV*�e�~/��yX\&����[���f��fQLLLL�Mr� mM� M��U�|����#O��8���~�E���{,ZbF�v���J�a��h9��6� )���v�X�b��w�!L�u?���Jn>]"��;���2���b�N�"����\#��w�:�M��?S��?�ɿl5��|�����.����cL��?b���D�E������E<�:��r{���,��H���50��^�XMC�����d�	�_#�����A���6a8r�Q��o�;ڒ�������l�ۆZ֖:p5^ȯ�\����Q8�az�0�+�c{m4��[æg�|W��JYx�M_�.�j����s .�h5XK{��&��!�A��l�{P�Q�'@D���ڟ�y��ّ��|������q��n�d���c���#����i��0�9ԅM��n�-NI:�d$I���ta��̽���$6�<F����@Ny&�=�D���f�������z\��'@�&�Bl�c�RC)�h�����;t4T��]�1 ��6�4 
���P%&5:�L�%x�٩}�UUltD�+]�&�9�7��	I��e���*g��kb�4�'�=N-_1�/�Iqt���)��B�7/[�T�/���N�����ҭ����or�u;�Hs��p1	���&��t[k���F���G?�K���Mi;u(2[<�zg�T+c���*�4�z���J���*TԶ_��Y���^��=��D��1@����NMK
V���]S���,u&��qÅ�^�4��m?M�5�չ����&�|��O�>@�r�����72��]k��y�#�����+�W���&.�O�����,C�8o�D��Y*A�ê>t�Y8G��^�B���N�Iؿ+pq*���Dw���2��aH�hhp��9�ξQE�����>�|B��>����>���[�ya�����;84�lM����$����J%}��$-
+Ga!_��@wI^��IVlF�$"W8�Q$�I�}��pJw�M!��?�YU]a�/������W_8��苙���ҰP�N�6/z�he�������(�*�%�"Nv��R�����@�&��݄��Q�Y}��.ܗIʌ0��}�����W�x����#o���X0-�>����F�~��;�8"P<KV�)�"I4E7	�
��+4�r �M���TBr5�g͎���U����Q�Y&�g�-�:�3�9���K�^�4,p"��*6�J2[�0��e""-�!&^�\��6�� �eb��r�Y@�\��l��C���}a5"�Z�ʎaE@�KL��M �������F�t2�:�pA{����pRI0�$�h$�Y �Kd�K쥮�������DI��AQN�T�v���ɜ�R��׀H�M��/�PW�זv��D�]�Ѱ��,�+���I��T��u�):��de=�h�H��}�(���qK�h�!���w)��Io�C����s#���q+l���$	�~@�0�r�nt��{O��6�S�L�^���"��<�Vj�����F���<|�^ry��p����|��P�0;�1��*6�]��Nl`���Ѐ2ҝ���L��'.��B���oo0�dk��l���+p��m��d|	�ߢ���n��-/����=����?���W�����O���!cn��1��~�nڰ[M�@ 6�<\l��U�~�ol�D-��cZ-?e(ANaŒ8G���w^nmK,?֨����z^/��V����.`���VZmǦ�Ă�k-�d��g"�uڄ�������jLH���� �<�|^W�~R���V|�H��+��)�8,L߫v����t�*�o90h���M�G�/nޣX�7�;'��n�{D�n���F����9�A���ōy�n剌������o��]���3�O]+S׺�U5����}��G���2·�n�н6�`F�o��4m6K�l�
U��	��!~����%C��L�@I0��ﴸ@�-4���l�WO�b�����>#�p1	l�7�T�aH߆Au��}0�	W�-���N��%SB]l��6].g�}o��j�+���5-�s���^,��,�"K��{ c,�Nb��[�y���+4��~���h��Ԋv���#[��D����21$�n����8c�5�Q�ѥ������Ui�U��]�����g��3�` ��bEt�u��I����鶱����j��r�뽲��l�]|ɸ�8��4&]�s��:����_���/�yT�;��x9��!�0ZK��b���/�'�pEma�܁�E���y��Q���4)�����'��`�S<!_K�r�iz��G#��d�j[�������XG�p��l��e��|-�.�a�>��4�Ð�vޝ��_�o�������f�z۲�	��@���J��Zˏ�ƛ-�S}����\O�)�^��ndM�&��&믺��� ���.`�nz2t=�+�E��e��n��[{=.���5�wd�3�K�������»�4H�ۮ�X���1�:5t. �Ǡ�ş�m5Lgԟ1��`Iк�����p>���x� ����G�����^���d3��zI� �)���x��*g(Ģ�� ��"��&k������􆾶2u;et_r���8�D{7Ϸtl|(6���0CU��$�X��qfj��B,Ds���{<�I|a���\(&���4�=�j&�֗^6b����v3��u=�o���#���]d�1�������e8�Fa _���/I�wO��8�S�ߺ��?�_�Ϫ�l��Y�à@�_�m�K?�y8��yd�}��`ID���*�ϗg����n���B�jΙ�bD�����Z��R���)�k�*4 ʹ�>Ë� �$�S�4���tCL�5���y�S���ƺʌ/ �db���j��u[:�#��{���������s�q�[��b����R�3���܍����" �	��{)8�bp����
nr���������l*�*�h��`�;~�nX��o�f*�����AI��Q����.�i9?���oK��7�O
�Lh$���/;��q������:���>����zpF8��=�xC��{���uu0p6�|JIIa]�S��9S��X����r����,�H�Eҭ��0���Y�=� ���`���B��82�����7��	�|n���{kT<�N��3��l�PŻc��'��p�Dd�7%P�,G��~o�/����7�t��C$��:i�K�;<��
s����cw��26�h�ӵ�ï^e�l�Q��)����xG%����^
׫+9��A����8X>РA��7��R��8�������1��䴖���B�7k�]�Ͷ�-Xc��V�`W����/\r���z.{�_jGC|1^0��y�����9�eD��${!�Kat?���׹PB��0Vz�����t3���LB�s6R����;���o�?$��[��T�h�������E�ea���L�����p�\*.ǉ#�a��VM*�34@d���
GE3�H�&�mk�G�sL1�M}���8��"��G@0������C�Rʋ�n�_轤���~x�s�a1^gꭾ�^9���f�U̅���K���D�L�ewI9�k�;�e.�~���9^��#t�]��0ŷ^�
��������K�/L�455m��K���2��ٽ�����>�"i�<��nd�A�r�p���YXƕ��z�N���:���TR������V�o�H��|����D!<��Т �p�}�	����M�4�^����V�>�ߟnl�����w���+��5	�FD<֫���ȗZ�˵2�/������7�,ty����������� �ǐ4�d������Xu��ٖcBFΦ4�p��W�d=�+��={�����R_a���[g,���L��Mжo��(�6&�#JƼ]����i���b���_��-������@a�"��r$՛�Q}Ѱ������V��/>"dڶ6V����f��d��`csZY�ŶrA��5����yt����&�!��c�N|*�)#E�~6Q-�2DI���ݛ��j5b܂��H�.��q�1gLR���0�;/���ɀL���"�?,c�W�|� j��b�%o���W<��?�:.q��=n�~�� c*�r�D�q,�_�u�V8UֿX!*�؄;�7������U!��l:r[`�V�C�l�o�)\�K)��0�v�wi�y��	�Yv�]�}y���i@��d*:�ʐI͕.sb�#�h���%X�B՘�O�Ӝ��:�����G�)�|1,'�U�8�����N��:Z�$�����*N�A�i�C���*�gZb���C���@4���

�}f"��<��]��{���ֵF_AC=�H��ߚ�*z��(���[m�m�C���������9��d|��}��v��`bη]�L8j�s?��uy������ר��Ld�3�X���|N}���ÝLw�������p��siA@4��{�g�H��M׵�,l.�N��Ơ��[�7]��=)Sʯ��D�]�J5z=#E���b9��r����<%fZ)dF`��d�Z�C{��{�m/�p7�H)y��N �uW:��1֞@)�٥��z�"�����7��\�_�3l��w��"t��dG��ZK|(R�N��%%!9r%PA����-��������6�к��h���E����]UV�o>2Af,��p���."#`h����l���"�y��@S��*j��<��e�)�8��&Ȕ/R�{���jCmOG����?
�II{_ܜk&(�k*������`jh�iXG���l,��M�w�$�O���o��ttx��u>'8�M�����~�/��[y�6��v�E���&��t�f�����9F/����Z��{kD�~�f�JJ%��!��f	��=U���q����Xr@=���+�9��\�U�Lq�٨/h�+�G�~S��%��$�����.~U���X��,�)Q��$��UV��5��[f���쮐�-Z)�d�I���P��M���r;s���lv:��F��9,V�j�ֻ��]�������{Nl�D7e��{=_�F�y�3Z��޺�2Ԯ��X�9%�xT�մ9��tj��vE�$��~�wBq�\,6�5x�a8+bw��y�*�_��<M�� �X,'s$���;N=$�A`�W!鯁md� W}k!�g���ʑ�U�
�eC5+.R�8����T�'��ð��5��}h~V[x&`�:�i��>��e	x?���~챹��3r�O�"i2���`d'ʈ�^^��������a�1���f�[������n�OV�lۇ�0$|�p���T��/<'͑�2�w���Onfi���[w�سJZcG^
�#��>^B��z��'^K5����לG�RB���;#��21���/I���j��F
�y��|_�������s'�k�{�6 �Q��Y(�H(`����,LZ��4��J�1��?����s�^Y�+=��G���D��m�у�Q�Z`N:�R�5[��	zaT��+T�2G�S�� X�E�#�8���Y*�J�ac�
����8���G�a|����y~��K���T%h�#Ho{�ER�|�w��bL/��������9��h�(f��%� ��	��9Ŗ?�������6�?��-s�L2�E��f�	>�r��1�p��A�� ���	�j��ʼ�Ȼd��p�>��\��ǈ^�\}e�A���g/��/��~~���f���]a�=�-���	�1�87�x��p�a�E��~F4q� ����+C��_���#/�3qD�ԁH^��L�C��s��>���.{O�}�[9mJ�/��f�z'��떬�.aR�eh�AOD��by��αyp��(��
�S���u����_���'�2]\����l�*�>o���{�B&�z�b�ΜeBn�{�l�o����+���#~N�р�9�7�Oq��#�cLK��`Ez�U
H���'�"y�JcddtT��{�4t����0���Ip�"��O�_�'S)Z	�=uf1D��.�+���)�r����
	w�G*����*g�T�tw��x\T�rG	�Q(6�$�m�
�|zeT�����C!����`_�0��pN$��"�@>O�>��T��屼���T̘e�~���&����袂횰�Swn� �����K{y�n�%tlK�U��n8�����u�^�<>�-0{�!�!Nn��+�{m�g�S&U���k'|�����m�!��\1:g�LC�I�����5��
O�X�w4�F7�Z�]�C�|�[�� >jp	��,�Ң��Dh>ѿy|�@�k_:�F�Oy/�^?����8]��><C�oA=?nQ�����}	j"4������z��>7�
�ys�Q�+�I{w�������n~��z�3�}�L���M!t��h.1�?��������ƿ�n�������]�p��X���W�H=����u��2U��<��u�3L��ks4V0���+���Ԛ�'��f����۴T���h<��[e�}�������p����Ȥ��6>W��C^��ԑ�^�`�p�Ç��c�,"�U����ް�С}�XчըT��B�s�;`������=�c��ӧ��zi'�0"h9f�;��{�L�6]�U�����}Œ����?������F�<���Q(�F_ߎ �
�o(�<��-�>[aXV=�34�p���BFͣ!��Rs�\o����Z��z��zR�q3�}˿[;�[��)�����k0�M�l҇A�����{����t�o��g�jH�����N�m�[xN\��f�-�_�w�]��A�WN*u���L�e��Ó�r"O�9�[K��y?�k�FjK!�g�ѿ}��-5Ԧ�_�p@�����ݭ�t}���!3�ϼvk��B�8��F������Gb����U�a���w�����رR��},��'8�{��P5#�ft���5�:9¾��x� ��x��P�\q�����"Z6��F�;�R��n���{0�57�$�Ӟr�+��4Ň�y��`�d4��� �D�4�L"jz�H\dus�߼�P�<
�c����D�6�=����<t�D�a��L*���x�2W_����J}u�Ο	kab����4b�R�{�����z�!���`�}�K���ߜ+�3qR��UmE����H�EZ@OӞOe󀽚�R�e{�0"2�ze��*�K"4�j��x��|����,��5x�8C��"�����Qnu�]���h&6�U��m�
<^�vn�U��6�Q5��������	�f����	}al#��QM����f����M�)-�&j�B<�P�=�,���G;{#��:�HO�;��"ϯ�=���Ѡ:����Cϙ��ُFaI�)��t��Ym�qj~<���{�ӽ��y3���B�p�mk�G%z.5����!=$$,b�-d��e�����,�G�?=����I*�*`�*�*����J� mUs�.�@��x.���63;7$
z��*^�)��65��Nl:�j��a��m��rPJ;�svɆ@�9��U#�C��X���ڢ�m�������zG�+(���G� :4zM/Z�q[�i�W(ɡ"�ߙa�B����g6ח���C���H���b,��X���$�:��~�`���)[0���}�IA�H�{�d�27�VyybYp�°�_K#G��9	X�4�n�b��vgj=�EAMy#![�~�ZV��HJ%	H�"���.FMHv��;=e'Nő@o�x4�"JI��Y[E����Rp�z�E��(���J���]��H��T�l��NC�ҊZ�}��o�U��t�j`�k���s/��1Nd{O"��弧�J�y���޾�>*�W0�n��Y[re:8J�i���Kۻ1nI�׫�v�S]��uR��Іղ������[[/��OEU��ʰ[�FƧ"�D��P���*s�D[��B�l���}	g8��&E��� F߬�S���} �9�U¤F�����d��"D6:.���	0]�<|q�NZW�8�:���@�Ӑ �>kҶ�I�!s�o�8�^E�}��T��V��N>D����l��%�%��\�SP�(��y"P����u��d �g�+��o��(��|��A��WV�ڰ᷃�H�#1�q�$*/�"&��߾��d�>� ex�w�+jm�V������h�s���S��Cb��"��aA�v�,�ʒ�&�Q�f�K�Z���r���eW,{[,�&� �L��tkts���u2�H�l��'a^"���O�e$bh�y��z����#�r���%v�����J�sLFC� �+�|��98(?H���u�\B.�����N���+1I��_��&��A�6R�K�ʨ}`i����d���N�"D�uL�2��023�Z�a�h���=�B�iF��������� �fy����l>�ro7����h�:O��}{���>�q,v'��F�t��p�������,Y:�!c��Yga�tM�~6Y{ڌdF��j?�������z`֒�s�n`�5j.G�"�G���@>�Ó��KF:�J��u�f4���ϡ�F�>�]�v���Š�8�#� u���\��჉��q_r,bD&�v&7��.6�� B���.�e�N���g�'�<� �;O��%�qL��⟞t�-9��=�+X�n��pI�'��"1+�!��RS �oy�	�k�ޝ�ߝFs)�f
x;eo�QWw��Bq����C�!��^d|��b�*6�T���]◦T�KG�\`A�_�d[������,*�ތ)��-̒f��n�n��$�L#T�,�H{CK�O�- �P5�iE`�ᬾ
�TP��O�������n���G�(��
qIǱ��H�wC��_�;ϐE�4		�;[�9�˝'���+[��x����Xf�D���y�5�Tc�GrX��a�d�ϑ1>�z8����#�rH����М=|�̦ˇ_���� ��9Jħټ~?�Ġq��3D�-�өfbp�}�A���:P��i�=�v��\	~\�����p7���b$:��d�[箷 �%ʐ�ܮ��3]0�K����H�ĕ}{��Ps�P�Kn��2?df1�3����шT��
Z��w|3L!�X u�7���x��e�EN��T��9�Ŵ����AH:		�Ce�F{�������;�<�A��J�v�Y�\���n�|�+�׺�}	�.!�̇ëἳ��.E0��$A���'�_Pa�2ܭg��?>�
�й�i�ڻY�X�42��&}3�VDZ11�h

K,�8�CE������~5�`:n�o�$Cdj�-���3�	�!���Ա�/�C�z�z(`�d8��(Ig%���@jm�U�a<�;�0` 3�Ϡ5>QT˷n�a#h�S'� �Y�(�I���xKF�ЪX.u��*����̤@$��+(�K� ܵ�:��S�f0��!��t��p&�\���8���-��[hB�^�n���dC�(�\M3��l�FX�\3 ,5���*�2�;Nj,���p�ߑ���?��}�;�缀�f��,&�"��5 �M<l[�pΣ���Xب����E5����u��GΝ$YL��6��@���W�ʍ���s$5��NP�eޏ�ȅ��Q���Ytϟ �HN���o�>'��<�i:���d��?u4�`u���ko#) Ϝ��ʨw�n��´	��������#����CB�ӳ$BpH��uPW�0<h��t"��­�����,ǒ=��Q'�Ht��ۀ
J %,pY´t	����p�0#L��x��3�c��g\�|U�V�	lV��)�WD���L}<��0��#FƟj�R%�e&XmH%��U~�����s��kk�p7�ª�B���7䂄���A��T7;��HO �$K�<�*��d az�=d��چ;�E@�Re��܄�ǺbE�`%%�s�Cf�;�- d�
��a��<��G�3��;	B�4�-D���	��j�rE�V��wY�������ѯWZ ��6$`��h!�K���y�,�*�#�F�q�Cf}��4����b����V�E���x�X��nH,!�#�{u���{:�`���������4G�*���ī�w(��*��=�Я/� 2,�Q�͞<ee���}��sX�|��/S�3˵{�#{S����N=k������� "X��@���M��UNB�f���&��F8r�"�a���N�x�1P�aR�٬�qY:PX�X�(�]��vZ4%�Рz�����1��#�Ư-�C�]a���L�1xa�Q�W6`n"9	�� {�r�p�l$7����C�'�n0�TH��JG|�c2Oj���2š���FG_#�����\�K���^����|�҄�7@��}��=V�|>���fnm�2S� ]uY S���=�9E�+W��mr,��M��r_)^$V�
:�ˁZ���+Aݓ��G���w'l�5�N��NG�Q$���(N�[g��Nҍ�����+H�+լ���t�rzh�7�7]�+�Hٚp�p�*;��9�Ɖ������Y�qG}N��`�heq�������vŭH��@�(!�[���N��U����Tf~1n��#��
���v*�~���kb?�n�#aC�MPh�i��ō��k%o�Σ�/ꂄ�FW(C��@��}�I+C��~�#ubAn����}**!>T�[=I��r�+��EI1��i�c��C��5�"G����D0�`݀	�'NN�.Ͽ�FbOQ�8��$9qpb���:z^�	Y,1=TJ�s�o�����pb�� u��?�v�5�����ٞ�B�����$���X;A8�A#"|n�j/�ʯ�Q�+�u	��T��Z照E�(��^�\P\>j��F�%� �0Jى8[8���D�����m��Byh���,�4x��E������Vm��>�H�3&ռ_78\�
��]����� ��&N�i�ۖ"*��>D^a n[�<��4P����:g\�0l'��)��]�f�� �l�c7�&�X���<F�<>����DRʂ5���VhiՅ�CuZ�O:��~$&:)N�nr�:Wյ�j����M2/���'Q̙em�0O$�'z"Y !\��4 Ǭ��'\A��㑱-��`G5�RS�2����[��,׃�L�W���U*��ۓK2� �]�Y��f�Θ���u��@���kʱB��WE�&��p̐hn2!DW�K-�WZ�H�k�u ��f�����w��6��O57�F/�e��"R �+��΀�j�]�&n�H@ Thf6NP�O�X��w�w�sJ��KYe����T'�"zNA"�k,-�6v`eƉ�ȁI�pQYb@"$�Ql�<�������]XXǒ>�v�V�����	�=M��#:��j	�i��i/�r$��5��Z�{��'�к��.�u�, �����x�ca6!�0:b��Q�,�.9�Ƽ��*{��n�5r��CF4K+W!�e��:�(Vo~[���X��x�~X&�*� =�VI���p�����AQ!�uL~?Vy��ƞvX�<�no�¨D����w�ΗPN\�ه -��HE?H}�s@�]|�0���3�A��H	�qߛP���(3�qi	�b�M��M��>�;�I�:����R\*�]�����2��|��l�~e��-#֩��Tu4e���8�J�xN��mGִq1��|q@�V�>�_�-)��˞D��8���P��4��,T��Oy�i���B���N��B����/
M�z8+Hy���#я_�Δz�}m4�����F3�]�Ʋ��E�VQ8�άn�\s��s���JF{��芬529G�E�`?{�Sa��`F�D!�Ѫ�����/ i&�,�ZU�v�<��f����S=9e��K6���_���4���I���	D(�
�&�Cu�IP�X����E���OSz��@� �\�
��-�ʔ�9A8�guT�)R`�R:*�^b$7�%fD�άԼ�?�.�0�(C�hA�Ϳ`���4I����ZŨN#"Ii�e�S���\�hq���<��7K�0*��-W�|�؀�k�����j3rIڐj/cG:xO�,��`,O�\��6��YU#�¯'=x�u�G�����q(�jhSBI�hJ�2(�:�+�r�$�@���8y��r��c����^��!kR���J�	S,��d�m���]�X�mD�b���#JL<E�B2�6ȴ�+8���/�$�DMd�I�񒬼d8Dph i�~�:�1���	�H��{�Y7*V��uI?�"u�B"��4h{n�����"� ���M����Ȅ@Fki��,��L�\�N,.�2�R��K��u��S��:[i�O�a���h�x�qH�Y� k{"��C\��&�-�^؇<���_p2�-*z(�}��':aJk$Y�}ή�A9�/Ԋ=%� ��c{ W �IJ �I��-���x�8C	�h����b����0���)z!?3�LO�����Fç��ˉ$N_�M=%���TTCu�$��B8
g�N8IWi�p��X����jy�@V��'� �8�L�ʁ��Iq�i���%��q�"B�E�씹]�T#��זXf�<���;cq2�VRLp3U!�EYCj)�U���K���a�X��[�#�)�\��E3��I )8����{��^Pf�1c]=}�ݹ(8g$�U�=� �������{�̮�+<��6T9���;*wmf�����?"6,aa�dk~����e�&C
>�0��Z���o�M�y�%�H�d���V�0A-�̹#C5I8���? m���23w����[go�=u�pc���~N���y�C)���M�������6~@�&��*�_��Љ�����̿bn�hK�M   p�P��_1�s&�*tAK��;�%xJo\Ir�s��n}6<ҧ�j������H�ԲK�(��k�����R�
X*�!�^˭)��@���ɸV���A�<	Q��c��j�B��G�={4,3��<��o�TΒ���~]���ַ��������� �89^XG(���:vNbb!ºr��Z���Pn}����w��xUz	j`D�T� �XQ"��T:�Y}�_�=D���&��޻��񳼪r�4so����zweuY��'�b醙j,dn�b�l��F��|��zZ	ъ��X��94����ɘj&����C�elRZ��ct�b��}�G���[O,_�!���,����p8+�峱1F�PJ�fJ��1�������Oe ֞9�� �|`//�Ѵ�9�Z�ʶ�hGU>��m+l�h	^����9�,=�aU��3��)�6d'4{��`$�ݎ���8wX��;{o�Y^,�����?�R){�He���WB��) ˵B�{����~M�Djk����ԗ"g;jL�V�z�֑�i#���'�[������u� 0-Aɑ+Hb��� ����ѳD�WWߩ~�J��S��gNMʼ*�xh���V�$��eH�[�`����%_X<�Q���1��ǝ��e�S��
���� ã����)�)�f�/�ή<���J���UHz���LBj�$8����xT��v�өf�^W���4�%��G�f����T\�2Ѓ����۹��$�/`�w'YN1ezE��{��QJ{����𓛔��-2d��bG�!%��V��'��c���-R��.�IۧwC��J[���?�� K�8"���(�T<�}!�)ؓL�=�_������I/�� ����2pt����*1PJN	G���Z�q�ߩ�kv�m�o����v�J+5kj[�AQ*	�X�Ҁ1�b�?6E��L��)ƌ`6c��D)<@�+(F����^U����"�7mZ���M�� n=}I['�
�d���B�N��>1����z�%W˱������V��Mc}�����67r�D^j?>:����9@�v-��bf���mj��՛��g�k�����@�$���ڑ��h���^i���X�<�r*i�5��"��M�w���+���*+�Ý���)@ێ�?����ea$3]zC�}���h	������0������k��ջ��� �D}�@]
Ji�
�G�y�m��8VZZ�
v�",�r�"d�u�Bu3 ]N��B@���U��p��� s*����l�>��WQgU^}ĖB�:�v�)���.��yW0�n7�)��E�� � 5@ʿ��4v`�����2���Dp����� ��F�IƧPX[I�����x�dl�lA�,��U�(«i����A���̳,+5��9dW
�E�P�EP�U�WĈ;D)��l,��nS�EX}��aJ�ZJ��Tc�����\K`�3>HD�@��E����Ɂ�^)D����x!Zm���q�𞝈r8 �����B�nP�Z����,�I"��� I���U��<���N!KqB���SY�������� @��6<���E�� ��^�����VxM@�G�jq��9�āW}�{���,Yf�Vd{4X]ь;"
T�\�(*E���?-�@�s~�,V�����,9mGAn&��(�UEIY�����Y�vfԒ4
�|��oƅ����eIb8H��¢	�p�0����`�ZqKEoiƴ(#�[�P��ϗ��e��A���.� dʲz�����፞�3�%G����r�gǬ��bh�yt8�R���F�V<�
�@���En���Hĳ0�����Ywb�b��GMn5p�RC��dd4�Y��$B��rq.|n�K�/�2�
�� �8Y5��"�lV��d��{�s�B�0x>�� C�,a��K���1����
�����E��IEH_Nzg���.����b7�5f|�?m�^��n�d��b����W��q�v�(�Ω���1�V(�^;Y;bccQ%�@�u�fW�T;�v~O!��*^�lD1���!�TJ�~�� ��摗uN9 �+
^)�-��B8�S��T�0�����8��6SU�;y芟5!�a؝.x��@S�QV��L�-"
�

Ir	؜�,E�\N�șR�^r���Q,֤�JJ%,Ui`�8���
fX=�.� VMi�Ç���w�m1h�aܰ����1���84QB�Chz�c��Ŵ���K�GBl|~�%�� wUv��7�_v`���3U� �a@��E�
��,4���)UY��[�%������%���w۟�S�F4��d�1��w/~>�°&!ʯ�)�y/��T�W$��!�;��l�����=����x#*D;p��l�{
�WLA��V<��N<vo\9*�������n'���m�j\)�D3�-�J�r�0fLu�C�euWM	q�D�B��Îe���t�M⾐s ���()B��_Ʌ�����`��u�~@v�p�F�8?���	����F��Jl��u_������ϻ�骓X�t�
7�M�iYb�?������a�kϠq2��$D�!��� �}�dWn���t���7�Ѩ�y����E;�y��EeK�"F����|&�N��'�2��0C��fY��B �P�����X�����jX��wtz�.8�砟���Q�6%(C�H�F�M��1"�ŅP����80��4|5�-N�00��5�v4�W�Zj+|�� ��}���Z�g������ı"	~���@$(��{�(^{�-Z��ؑ�����K$���3d�cd����6#����i��倡/<��7CF|��X4m�Þ�A�xb�WP�D���O�6h|+��W(�p�՗�⦚@�^�#�H��CŊNp�
�'�%�x�ջ�y/��;+� �ŏ����V��	�!W�A�D'>x;����a�����-&VI�S[%v��b�b6� �,�.aE>Kgc�,c��A�_��o��8���K8��,�O���CX>�N����1	I�����������l�j���д��7ǰৃ��*�X �6IE���x�#��>s/�+�jg���شu?gb�,x�n��q���
bB-���D�1��Ag|�u:f~���6�˝+����ps�
��A��1�B-L|�l�y��	��#F.D�\�A0�������hy0x�R��p�Y�:��l$�|���{�ɗ�h�AԬV	s�ނ�Na��D�D���[�)(�e�II�X�p�ˋ�T�I1�s�B��m��,LO1�m��Wy$���ހ�cּťf���.��d�h3�q�DMg�J��N3���B�=���"��Cg� Uv�A��q/݅� P�$8�X0a�/ظ�(��ZX+�Ч���vR�ɦ)�/4��y*w��O��~���20k�T����6��H�y�� � o���G>ޜ�5�5o��g�`��?�L;ܼNA�uQ�tޙ�֦y`�;�Ψ��(;_~�	�v�+>��g�ʨ�Q5	��\���Y	7��wc�̧���6��\����~�;mʅu�GdN!r
��*�����e��ja�;�Κ9�*�"�f{
��L�OC�|����g��w�|sؽW̕�%�f�hz3�o�f�"��Ҋ��:Q�H�Xr)�E�X>�$��S�!��u��T0aP#��t?��v5���3a�a`�K�UD�_�hs��5���H
��,�ۇD!���y<=�g�~9�.�ۛ��E���' �Ն3g2�v2�>�Ʒ7��N���Ե��ޕ+�G�
���M7e5���Mj.?mZ4Ľw�@�x�D�ikp #��tB�$�g��V��^��
�r����[��Q/^���I���������Q
�x���P<���STMoVә݁��~����D3;M	>���:� D]a=G��L�&����o�r���`~<K���-�|7Hc�L,�W�k�`�#
���A�M��qmp����o`�������8�)>\r�mގ�BZ�����������-G��*2����>�t�����0���r.�!���kÞ��{�v�>��V�t��We@�B�T�F]�D�֩�W���7�bO����+p}���5�����2�(X�~�"�Џ�n����S�u��Wf���=��7��}�3�Z�U��)D�X�%����M�xuc}�? ��o��>�qp:y���)�JYZ".�j�X�~0�μb�ӹ0Av<�6Xc�S<9�V��בD=��P8}ʨ{��z���c�r%��2��f{F��Q ��Ϻ�ؘ�O���a����1��� ��q[��i��?=�����dx�{�oEy��>�Wۍ��  �D�5zMrb,�'1���!��bb,`T��(��Q��J�}o�m�5�f����f1�lr���{��/?vYk��{�Sښp��Ǡ[W��ѯ��աP�H$��=PC���\`!�t�2�b̩G��6�+_��uM�z퉨��z�ch�I4�X��-z�ի���sg��e�������b��f�Y�q����n}7�ѬőN7�[}5�LNf���d���٘�����3zcƓ�1��9��H�����8�'&�p�;��"�}���w���,��s���و�yD��lT�
 Huv
A�qw$m��{(dp��mb�)�V+J���9l���g&�܁����RVo�ō��"]KS`����pbpCj�h0ۖ��~�ukC\pǟ���Ǟ�\}����u���"�t���ڽ�\8�	�>�U$�	���������c�1�� �M�vܾ��Y�_>�M���>�L��� ᷼��2�2��ѳ��Z�i�/�-¡������'~�W��k�
خ:����%���X�`Z�w�Ǳ���}/���]�Љ�s����Of����������|�5�/�L;�j�����`�7i���f�8D�)�k7��+�}�1*bs�Vj>%ĢP��#S��'	XKo��afM���ч�{�ɟ�_�^�#h߷��A���CJqF1�Je��(�Zгk0ᢃ�ry�_�0m����G�\����S��bA��w$v����N39�j��f7`�I����ѵ�Ud}`}+�����ݹ˰^�AU2�[���p�	?�N;*��������}
�]�~;����{	���mo����c�	;�Gf�/��G�����L�:��ޛ�O��v��S͆�p�ч��ú�*4n ���	��fu7�;ءg~}t?<��\|�,#�	a9/�	�.�궫�}#\A�`���B�sS�E[�& �H���JIP�m���`l�v߸M�z��^��-%
$j-�R~{#�����:#W���,�N99�M^s��$�V~��c�S�(����Ba�n9�B!��]%����L��B��j�Վ�ֶFxe6+� ��Ч_����-L�d��e8��ݽ+��V��oB}C'�c	��[��Z�e�䠐P��A�J�V�mCn�h�&���_��J����:\e��",听�C{فG�	�w,Q PmG��E���A��p��X"H��E#z�J ҜiT���d���ɷ�:��ߝ��wf���mM��H��ٔ�*�3E��@�z/�4�vL�ep#�74��H�P�\�^��"րnZ(�J�c����h!�%O����8�b	�W���V�%�h��ajUx�e�ښb���2m>���t3&���Dܹҏ���X�d;��x9�c&JtR��(����F�YJK�P�G:��lG��!���x�$�fR�|�ݲ���	��	����Qj�p����'��L-E�dmR�$U�n��1���1&�ҁ���>���9�����y�d��$-�N�+'acȴt��dWA�-�mn����
3���G6�!�Ƅ��#l(�uUӰ'ס�x��v�|*|�Y�ܶQ�J�S�6�@��]O�4x��\�\l���<�I�7��䁍�z�dP`K��""�<Kn<�<bF�ؒ���U:���(�]L��T*�#�E�"�� �]S^�	�� �u<(� 33e�Q*�?C�1Q�d[M�s���!�������7�CH~��e"��7آ	-����W�oƶI�-��!��u��x>�)�f����6TgMԷ�	9I�o���p=f� It���/�1��K�G�[3\yR��!�nh0��O~��9��Z䒭X,J��m0����.�E�%�տ����!,g�f��R�@��-@gG�qHt���'�uHPY'��Qd�P���E�;���|^f�cJj%�M��tb��N�,��QN�^�ȖCՂF�1�kW���c|��h�j�(R���K%��ǶL�t״b(]xAI���'���Ϫ��L�$�.�\oe1Z�IV@Wz�P��u�✘|�i(���h+�$C9�	![y��W��1C�AQX~Y�wT[�ZaHU�DL�e'��t����d�"D@6>Qi$�9���Ǫ7�D2[�Q"��V"�A�U2��䁂��#V����y
�<	�0p��3�U0c�eP	 ��ј�R!/*ER\:@�'˂K{�h+�u������|f&�|ɖk�)�>�_C/������!���	S�±SR"��v)'�1W�c�O&�-����8�����)�D&f_6�B�3����(���#H�g\1�q;�4e4��T !z\�.ȶ��ݾ��:L�$�/R�N�W*"��(�����tH\���ֶP��4D�e��W��u(�T��ĉ%%��R �%��c��]Au�A"��b�E�ku�ĥ
ZK�����\}+�C$j�F�at ;Y�t��/���FC�����nG�ן�~���Q�Z�+��. ��z b��5;���Ү*>�~A�V]?�=IU1�s\d�H�e���e�2���B�g�@	����6����L��;�z�=�tx������.���%[ذu9rm+�Y�����(R=?��J�Z���1��}7�2Pg�%C�l����X��2�f�`��T��mҷ%D�+�E���kuEu׾(���ld��I	�-�L��.A�V؊��M5��{������P0�P�g����ڜ9Њ�Q��,�
ꊆ(�_`�`����m��&��D��bB����R���>\h�*l��P�{ �e�%@Ls��rff��/�EˬH���ƀ(N�DgY�`x����]8=�����Ku�G�9W�e���p��b+��J����1P΋X�D��=����s�bS��?O���@1�������2�����S��/ zFv7`w�@c����z����8��?�4�1�W���G	�s�E�O!Ձ���$Y��I���f�E!�p��Opc���Q(�b�LԘEH%9J��1c|zǿ!cXAU�&|6����cp��=�d��|�vL1�\W���$V�g1v�8�<���?�F���ܷ�P��<�|�ƣ�g�8%�(f9єU|S8�=ޞw��{s�ԋ�q�Y�b]P���!08����8:mh�x���q�Ǡ�*�|�m%S���W��e#!�SO?�O�n�.GCeyƓp핑r$�"��,v����G�+�����{�$z=pᖋ0l���'^�����Q�E�Q��fɑ\��������gb�������
��I���S%-�G#k�����%M�v�c����T�� 4���cף)B�JIԇ-�=����5�*%��h-�u�E�`�Iا�g���b��y��ȼ�I���/�N��A��P�네3�����������1��?�� jw)�(k��m��%�$^�KL��"{��)�,��z��~�~V�}z9M8﷿��0bP��,�T�B�d&�1��'��7-���+����Z��.٤�N/�ӗ�Ð�&��ݱ�9��C�84NwI �4�\WP�0�x�Y��4���9��i>0��5u�$^Z>k^y��]/L�
�U�]���CA���j|2n�n*���.��H����2��C�ƽU��i�!l&#s��K�<ߚ���s}y5޻uι�D�kI��ܒ~ԨL813m�/�!�<�*�=a,�>��Df��������ܗ����0��?������JA554���o�|�<��d:������mH����t
۰���7��O��� �BG��XX��bP���G���K��㗗b}P'��m��˷�������0(���c����������%'�(=�׏���=�qH$�N��P4ѫ�����������a�%�����A��(��TU>�|>n��A�7�����#ű)]�(橮$��-iW?�cx��ؕlm`P���	W��O�A�v�
[�8�}��b��n��n�N=�bl�a���@ul��ٝ��r3
_��E3�Ľ���sr�^!�G�w��C�������ć^��LC#:��'�&�Ð�7�?V̺=�\z�)(�R�G�l��lT��-<��ۘ��~z�zW�%�a(PL��b�[�`P|.<�h��,J�{��x(�B�(�D�������c���E:H�d�����!j�,r�����'�����Y٥2�i$( k)�Y5�v��.ĵ�c�K�Z�f��y��F�
�CK2�nz��Ç.���}+F��U�o0{�8�̟���n�R��J0d�� _,�w#��N'�n�]���/���o=����.����U`�&&
ӌ�+���G�c�3��Yw�I�8�F2։K`�Κ�[�Əu�O9^�����nR�������k�t�p	��C��rXF������=�]��8�!Α��L�GG��G���'I\z����W%��Yh�(0�Y�	nM�An��X��$<0c<�0#T���^�v��̆i��}�?����h:�esVS��9ͷ�C7<t���;:[#���训�[�/A�6zVs���8��#��T�$�d\�m��9+����a��[�&8̒�@�'�d��g�c�돠W�ZQ���O����a���L�T��M�7�1�tkD��*�0c4|���h��%���E�n�-�uM����$%��A����v'��Xl(שVT�(߅��]w1���W����@)��g9P�!+.�Xt]l4�6]    IDATZ�G���=�d������	�*0���#��N��$!8w�]" 0��eőI�֬�2����"�r�g¢=�f��Q��#2�n�|�@���N�2��倷��ӈ8GC9"���'���7ջ��(������>���� �44��$c0�G�Mōl��z�����J�1����)��7�OF�{��K�
�*oL�����
)��j���������(��B�́[���/_�抗p����e�2��t�n�$�NSs
�W�ÂFk��߯G"�Q���-�d`�m������Nئ��BlM 5�RZ=p�$�����Y�A܇l� �=�Jl. %��g?W*r���#2Sƍ�2�ok�:�RcL��Y
������P�{u�D�^�\@��2u���y��w�ᱏW*;�$qL�����}/B�d5�$���u]��P�6,}{Z?z��6(�]`(�;Ճ7�1���h��Q�Ff���Z�c�;c'�K��!�٪(d���1[pc�����o���6�S.C[�V�y`�-�-x������
Ze�*�@^�� =��ɮ��kZp�3��ЩhM��zEށ�HW<X�>[S�B2��!c�K�A�o��Eӊ�� �E�/���t=n4�|�|5�C]�@mЪ2�_���xE�>c�I`�.�V/����tc`p���uT��X��T9JPhS�+Jn3d�o��p�a�?���Z�h�Dƽ���Z�a��b��|�8��\��v��.r#�IUk�������C�þ�C�슂�XJ,�J�+X��x��?�����f�!��F�k�1|�]x��T��pK�:�)_)V7k�.�:̾��ck����G�Qbjō�sN$%}tbYj/O�	�l��$1� �Wc���W��lW[T����Ӓ1����(ql��0m�?̞�k�#hһ�d�Na�Д��1mt�rX��$���� �m�K=u7A�T`��AWs�C���c$0Ȱ־؆%c�k:�H��'$AL.-�?�dZ��+K�/{<����U���E8p�uh��Q�و⁰]�`nn�_��������7�U3g
�W�0�V.o���ߏ�gޏb��pEԅŪjUU��L����%Ό��_�Y�������F��hYf��c_�b�fg���eH�t |���\�X��3��KX����%RXE��'��(�U���$�%�e��֎%o݃���_6Z�o)c��<J��NR'>Da�:������-6�O={)ӤӵHʜg�{�rM��xa�R<��2|�x�h�ȋ|�rT��@������Ϸ������\ps?�M�!V�FkW�1�ҩt�d�v 9z"��Y�$,����l�J:[C8����������|�΃�=�.<� 	���M�h���!�!����K��c+qȹ�Ь�6v[��6�翈�/܊�R���U���I��r ���&��L��
C�ƣZ�ہQ)>�gq��}��{�}\\��#z*0��c�o�c�D'���*��V�]���7���'W�a�eW�)c2ǨC�
��o�\�����G�dZk$$0�����}�Ԯp�}*cc`�(��O�1�&|8�5����'��Y`l�^!v��o��Q�Q}��c�;ӱK�s?y�L.��SGh%0���3�%0z���=�Dʄ�oC2F�(QNӢ�-���}����r~�!d�v���^�"5A��*��%�����*cl)0��І%o�������of=�]b���S��S��.���&Vn���-#�g�X���^�μ�F�ZLىs���$;�%,z�VL����ƈ�π�-�-����vu#.���{xc`���f<�X\	.�v�0|[`�;���E�?��x��r�hp���ܩ������Ģj�x�k<�\#�=��#�(Q`]���7����W�A�ƨ����/��ƚ��(r�ChO@��*���/+̐�f�(08����qS���?[|n���]"-�h�!����(����ͬ�%1眰?b�n�$ ���R���T��*O����ԂCϾ{��0�!���ƌq����I`DXN����5\|�r�	�"��� �U����c����jծ�WG��q�TsW���x�Q�nǏA͎Rn]�Ս6!d%����G��g����sc�*����yMܮFʽ�I4�����7�`���C���f��l\.�L8 �0w>�~9�A'AZ�vՐ�j�YƂ����g�boh��"x��U5�㢫H�.k�x���x��=�FlM��Kl�.]I-T`,~~n��<���;�!s	�j�F����hn*���f [����*��H��H�[�0�%wt0clu`���u˥���׮��
�D�@i���Φ
�@����	c�;��D��Q&G�z�Da���������̀p8�D���� �L����P���^8`��X��;aœ�������q�0�E����J5��X*:)�X(�}�tv��H�]a�`�� +�8u�,���ͺ(m��nQ�{8	"A��ϙ[9Qt=��8=!:�$o3؜@C����YX����(T f��m:x=��*��C�`uƐKF��[��U����&�Lc����P���1<�!���|�yԖV��)�����Ñ��Ќ�4�0D�����}�DJ1�`�̳Ǣ��Q��"<V�q��d>���.���OM��i7�*ge�,�]�����cq���LL������bu��0�sՈ�4b�<"�6`��5}�+Ǝ���%]�D%���2�MA4���<�����Ϯ�t�d�Ő/;���JҘ���(��Pn�n[���^@X���iZ�(�C�z'`�ð���G:��lR�}�cA�xi���c���&�8�%J|��.Ǽ�1X�eW$,�FW�>�N�]	Q�X_P,(����C����FW����/��'���iׇ�,S����1�D!���:�3�^��'\���{��ɹ,&wT�R�x+��WON���7���&Q�m|�Es������[31m�+8l��X�s���+�	��t�f��wr�?��7ހ�����7��6��$P٘��s�˜����[�5�����<�q�bէ/!\�
���2.��8
W[e��{ �F��W?���b�翇"���)nw	��׌`�{�������"�N����^�!���������и�<���06X=�JMXW�*2��i���d�E��[�]%����s-~w���>��0�O�N�-Sp��G^	?DU���`�IW��;�:���g���!��ފ���wb��7
�U��h2P	7��ƛo���z��=��t����Y6���d:�����B��R����:�nM�|Y��1L�Y��4��^��F�b�������ki4��+�_<�i׏j �°�
�Vf@9ЌLC�$�>�&^��{��9(�c�-M��@��_��z�VL��F$��rW"Z>r"I�$�S@��͝����C.{��9��_!��5�%�a�n(.���YcL��#r�[�J�x��
sf܌���$O'1���Җ��%��ō 邇sG^��']��n0�<i�-�Z�Q����]�}�nL�~���hW�5*�c���)+���x=��>���]ap�	��j��Q�7���h]��p�h$l�|^p����@��`Oa"``<�>X����^�f�q�\� �]#��x���9o�<�\{�Ŝ�tX1d�98���� �g������
{��TC�E�s%�"��E�1wL�Ն+�!&��`��D}J+-`���q��ǰ��I�$���hZ�0�Wծ�����gv�͗oY�sk�:�NF>��z��ȁ8���D�F7
��ȵ-�����$�<�Jl�eH���+��LS.\��
2(�x�w30�c��K��z��2�$*q�iZxc�'x�Y8�;�����?d��P����P���/x7����F�����`ծ�M�l���䳘��Z�s��h	����h��^��z��(~����r�6�P"�1���J98Ҷ�¾��ԛxc���q6�<e+!�L�N��O�[��>:�M�*��R�n�w����Z���/>����u�DdR��Xr�P�&�3c`H�U��]I4��Q�52��׺M��;��z�B�{��r�>��
�F�1�k��/F����(��7����OF;r+>��Oލߏ�f9#P>���� 
1z=��{}�'��9�;���e��� �8t��zvγhZ�.��L� �`(-�1p�LN�3�^���Vf1��ñ���G$��47���_�	w�L\s���͍�M��x2&�~>��GJ#q'	����xk~��rZ�*xvJ�	nbƬ
3pW���L���nAJ��&��h\��|���O>��w=�C/���ZvJ
Ve[�D�,,�EeC��H|�ٻƏ�ѹg������?P�ٚ� ��m�g�4/�P��\�7��*��h�����w�����"����5��kHy�W~��OL�,@9A�0�s�����
�ͦt�{�~9�5ZY���PS�;�e�9����y�)�
�z\�i*쳍>W��ό������3�E�������O��Âw_D~�Ӏ������Y#�+�wJ>k�w���Yhu�(�D��`��D�5_�GJ,>�AQ�d�.�]�l�M�����7!��A�>?$mG���䐋-�V���W�(��_�PfI1�*1']5"�Q �ݪ�!w�SP�����p�6X�Cw�$C+�JǮD�v��m��I&�Id�:x�S#=O�O��LCa���3(�����Př:��� $7��L:-w�'��������H��ڡ��dh&��� �K�X�{ ���q� cA�A��,�X��6Ӣ��+߈r�(礫���RS���&
�r��%��V�u������T8��3�>F�Av%�]ݚ�PMlK��s\�E�vQq��"G4?�c��Z93%�����dh�	�D:�t!��%�>DBHɂ��Z
�h,�(g����F�r�f4Zbmn�'{J\��4	�ȅ��
�h9+%�9&��X�j�S�G�\D�C�D�R�VY��5���j�*�[�(MPC�5��,^U1�4�*���G�Q��5=JF��O��K���HoDv����F����N�����KYT)Zn��ۡ��QZ���O��dq�)T�@���``�W�GR�\`ZaF�!'KD2�7�!��vI�óU<\I�*?4:-Ẁ%EYC��5��*Spefǉ!� �d
�� s��nW���Vv&JF��7C��L��>8�si���wM�2�4آ����
��+�X4VG&�Id�DEHyK��B_�B�b�A�N�&|<���qc�lή�a�8N��LJ�GE֖�O8J∁$fp*�q��񆋰�����	�;(F�h����E�1A?�5��Qe&U�(?CYw30x+6mJ���r+��H9Ϡ���d��qE��d@�x�"'�x�����H�Ӕh
	?�A�h�G?V>,q���SX�>W0��uTΚ�<�"j���=l�"J1�;"Pi��cgS`��K��e�q�O�9�w����羇r��^�p���E���+�n��7F��se,���QN�܍��<�B�r� ଟ�H\�g��cD�YX���� �y3U`��T�/t��&�b�RA+�e�j����<���Zo���yLX�|<.D[e�d�<�|���`�̈M�q�������J�F�|VTT�#Z���f��k,�~����U�%�kb���_��F�0�Y�D�v'�:Jd���?0$��jW���RW��M�'ʶ|���QGwm'���L))FUᤊS>J�J�C9�#�J��O�T]��U}Q+N��h��Ŧ��V���C*GG�1(���a�5��H��V��,<�� r��p�$yE�"_�~��<�f/Z�c_�1R	�cS��UQ-���QD}~n����/T楊�P��7�j5_��m�*>͍��%0�]��0o�|*K�
kL.Nt!7��Q�D\L�F��H-��,�<~ʏ����0��i���>E�x��,R�Qe����Ճ�o��0��]P*�D��v�v�8:�虁�T&=<�:\I&(}�YI%}Nf
�xx|H���[&��F+1:�YC*�Q�I�-�3k ��{��M���T���Mq7EƔ��*G�a�{D�I�ԋ�Ht�5�>�L��2~�k�i�fy���_���$z� Fda%$ y��gy�� WD@9R"־ �&�|�����B.x�RE���UlO�K��At�J9e>i��������.���{�*y�6�n\Ή�w���@��ZW܊����}��V�P}$�I^f&Փ�5��B6�Fbv$�������fS�j,�U sr��ḷ@�����"e�����ˢS�g�L�U�*���Z�!hפ���x�'���o"�m�#	��ƿ���N�W7����sjE�&�6�+ ��_Ԏ�8�����eJ��w!�	Ӷ�泈9Ԩ����F����rY%���!G��g.<7�H>�eU��p�u���:M��d�Q����S�CPwӎǐ)����e����ԓĖ��\����J�@��N"��Fw�جZc��0�(����%�^�Ϩے���Q�]�Q�ߩ ��3T'�^�����p��ZLJ�D�+����~��ˎ� Gn���:z	E������)�;��<0�4"����e�w��=�PB])�����/�p�У�gY	����ؘ+�q��P#E'���E*���2��)����Z?�[1�G�"�T��ȕJ(���;�QA���$� vٓ��O���,��*�b�Y������ి�WZ�ddN���rQ���ř��9Q��/X�Yp��y��ٕZf������k�����W
08�|)�):P<�|T�.�&l~��e,����}�y�:t�ɟw c�$�I���r��(zE��h��PcI��>)�Y ��E8�����l�[�s#6��b>+j8��EN�"pRhn/"��H�yT[�ީ�Y�n�RI�VR���� ��D�4��"h]���!i���e_d�S19��t�o%�C=z��rU�0Ljp� �����D|U�ln� �K�А��r������m�U��j������P����t+F�(q�e��P��ކOo?==����)�30�L�q�ЋT`�G��,ʬ���վeb������m�ߦ~����5��D��jt�H��֮Z�uO�n������) Ā ��/��^�\��;��mR3p�W���� ����ߧ�~���g����? ^���m	��~:����g'���=��hhk�@=�a���3b�Ӊ��bI����{�V�dQ(f�b�����؄��
�$ߑ?W6V;���S>����IU��to|�2 �!t�<ЬYX�q�������a�n�h�s�8��-�ŷ���wJ`���<�̟�}��?�;�E\s�0�n�I4���E�[����?c82f-��.C�����᧣*��!�=����m����Ћ�AZ�F,,�����нk�,�x\P��ؒ�0��I���@�'bz�O']�a瞈���F�Ǜ@�=��6�K�n�Cp�1Hl��}GIOS����X�(ss�|ci�r�Hؾ���~�Ѯ���Yx�F^ ��TZ�ʤwk����r:.��P󞲡8V&*�]TQ�4\ɦ�N}ae�0kҘ�)��w��n!0=r���7F,Z�t���q|�.~M�&c�u� ȳk�P`�Ӱ��9��F_�Ç_�l�;��E�;�q��Q*)�5�I���_���u9\5�&0�jd���i|t�Y���PW�I::'��J���>���$h�,���]�\w�Ht��M�b�]�_b��%�c�� �Ͼ�Z5���^JY�F��m����o<�`��$������b.�,�D��ǯ�АB3*Z��T��D���Qc\v-���<�Ja��F��^����)�H _n    IDAT��r`L��5���>A2�Fw*��qѡ4�,¦�X��͘���ÆǳMv:V�p��q8�?�9�-K���`�b2�v�w�"eؖ�ōy���Sq��k��o@����[~��:]z�Tn��}�]Ӏߎ��G��t��Pk���� C@��q���SC� di�(]�����.����D�Aڬ���E~ ��5���%T�!�~�6r+���N{��������R�t)�#E���������V�r!Tn��a5_2�ć@=M�\u�����-���F����愑�S�{�g�����.�7md��Hī��K��c���q����2� N��� vqc��D2�hKl��_�p��I��9���N,��0e�p�Tr�MXo�@�܌�������.]�t3��Db�,�4g��=~<���V����N�M�G�.�jmz�5�� ��8{�x:�7(��mV'��!�r¶��J
��KRp�9|3�֭��CQ"�?g7#�P����;	�������h��uߴ�Wˍ��7����۰��u(��%> l�"��D��a��/��g��]�O?f���>i�w%��y���G]��!�!��'5�$P�*���UBn�L�|�6<x��02=A���t��l��އ�-�Ѽ�+�߹��*O)�8+U�|����a�~�$6��	��[���ᦫ���[7�+(�H��bX1\x���w��ж��b��y6n�r(���	ߧ1�����A1���+nĮ�ׯ���j�2�L8�kg"�5U(b�ϡв;>.�n���Y�W��+���X<���+�Ҏ�,�Xl��L��r���"�Y�f��?F�b�YW2l����n���-v%*0���!N�zԉ���q]"A��0���oc��ɸ��+��-]�h�h)��e�q��p���b�����c�_oÌG���#�K%MGm"�EkҸ��;p�W�X�z~>��t�t݅���C2'��o���bI�2l�����:��bָ���G��s��� ��I�z�F\�}~zܮ��uF.�e6!$��إ5�c��O!�Ҍ��OKD��h�(��j�*���\���d
���o���h��� Q�r����2w&�\�O+�O�Ƞ}��h��)�I��w�<�}��1z���.>�}��]��z�A$��q�H�W��Ϟ�.*2J���N�c<�i�c�U7��F���B�j)>Ǐ��,Kj�`�r	�(����f�q�yi�q����O#ѩKW��p���i� �sɕr��ﳏ�-�<�R�r�p��7.#���������O|�Q0z�\�rNg���'��U�6�a��#�܂���	\����Z�݋�W�[�"��ʪ��q+�cK��nį�*"�c�U�SE��V8�72Ȭ���9�c��k7|�?���I���rƘ��މFԋ�,�Ǧ�"�r�x��JM�.��#��[P�P,p���C[��ܯ��?%��r�V|��A�vqF��[HB|��$v�y$7�(|��k�uie���+kh��;}���;�K������y��CUu��Q�.�:C<��y�=���Z]_R�������wV��'̰��ȥS]����E�����%�F��j,�\"��R�������޶�����T�&E�BU�wZ��d`�H��ȭ~k�|�A�ƉM��m��Ʊ�w�	�;�1�~75r:�|������ yq�!��2c�+^X��S� ��a`O��� ����^�h@f���*rT�*�����������Wym��y�op����g��9�Y��O��M:��[�Z���E�^��lK�r
z�,��U�R䏋�����Q��i��ŕt���
�韼8W�Qo@$u����|���H�iV����nD���ĳ�&�u���{�{��3G���>L�F���y|���(~�*Pj�11��!��Ӱi_�`#��T���-�~$��L8�ݨ�Z�ԱPR���M�'��'�X��^v���d_��~������y2�R�sz��w<���*4y5HF�'ї�3c00x����g(j��J`Tgj$��Ѱٗo�P��e��E����^S�6z�S0����QQ��MT�mȯ~Ec�97#n���1��1e�#�9���O��A��ڰ+ߞ�?[U,Tn�T=j��p��1Me�
Eo�����4��=A��Wc��z�	eSs$�V,�D�5V󏲌���B�ΫG�lu�������5?G�
:g��n:��Gl
��<���D_G}؎��@������V�By?ɵvEZR�6��Q[l�eC�yM�Q;r�ȕ�����A2�����&�FJ�^Ɗ/?��a��1C̾�ܶ;o}����E�����!QX���ߏ5��EP���iM��$�@��ʲ�B*7K	H�/b�*�XL���h���h-�D�1sk+.F�d�O�	������E�1�����U�4A����@��� �_�ɒ��A�09J*�d����5��ϐ�E5�ڕT��Y9"3G*Ҳ��M7D��:rR�����_�
C��b�QGö��$r<ʨF��D�I7=���hcq��j��ȶ���ӑ�[P\�*V~�)vv�pwgO�6��Qm�]�z�?;����s�9J�%袷c��w������J�<*�Y�������Xe���:z��#�n��Q2Q��+�o}��n�6
�Ejn������=O�f��@����y�}������������<
%t��a�p���"7�j|^q�L	��M�TA��(�@(��O�Q,{����d09�Y�T�������!(;ΐ+�2}1���.j�k�Q*����]Wl?.�X+;J�Q�GU��.i�"��-���s�~�8�u�(�)�F��vu�O�쬋�v�᷋!
U��X��d4}� _Ā~c���&����6\Q`D ���S�CJUc�������lt�AfxCd���lW��d�=���D w�C��r�(�[ø@�C%�O{��Eo܄���hZ�ɺ8R5�ZĬ�̅ׯ@�ϡK���)heq-@�m��M�Wա�~�~��W."nSۣ���Ĝ�VJ���!�������wb�"a�!��]	��î��������#�=�-0: ZDj&���.��$� LG��Am*���q�b�N]�u�V!$.��G6ׂ�_D�>}Pv������epةK7؉*�3��H!�H+�ǆ�b'KvB5�g��e̱���H`�}�Ň�s�o���Q��|[`t<c���bNc�%e�+-&Qd6t��$@�Z��������%�;%�HQ�\C�i���	͙ft���U-{�L����X5R��a�q�n ǈڬض��ص=`�ꐰ���,il��2ƶ����EdbQ�J,#0���D��Cw������"��:��>GU�ӱ�f�R�.Q�9��T�����k_J<��g�y�X��ֵrĕ2^�K<U��E�L9'lE`�O�e�!g�~ʗ�2��Vc��͔9��3�	����ۑ͵�h�[�ż7���K�h\���z����~{b�;!,瑬������,�[odJ@]�t0�^��b��ڶe�'�5�K�2�$ I[� � ]�t���X`L���qC/���m5FGj��<�E�̒#@!�Ќ\a�����n@��yX7�E��i��ð��H8:���!t��HR RH��X�f-&M��Oޞ�Ԡ�ѵ��j5XղN�
U��H�k�20ȋX����-0Tq�q��NWB7���(#�s��mhA3��%�
��ڴޒ/D���}1��Y��t�2��k�����r��q7�/~Hv�vA��.Ы�Qݝ;���Ȓs
>�f%�q����e�m�gǋO.����Lő˷�n��Bz����n��/�Ev���i���'�
z�ҥO?���Ԇ6<�G2a�-�ʮ��;'ބ��yI��v�%�k֖�������+Jb�ǀ�ʐ�FB��hJH��]|n��{��� ���|#�$��!��)�cݢYh�`�;dw|��,����pvۡ�?�ڮp�	����T�
�n��?�$vؾR�:|>ov�7�7����a��G�h�@10�1������Q񹱘�B`�5~���uҜm���T|���	
�X�~B��TM
u5lw=�~�~@[#׎�{�C*Y��m/u,Y�5vݥ?�|��;�X,�;n��=�,RH�-��yTW�b��ň�vG[����T�G��i}�X-��pI�)nޕ(��p�o��]��G�F��j�ge^�Ѻ�t�3�塃1�曰]����j`��siT�m̝?��&M��rp�mwcƣO���3�V�/+ee��_�#~zjz����?�����������I`P��(|%I��%0��ķ��ಋ�������V��^�����57��Q��in��ӧ��v���HC�|�,�f.~pȁ�a���6�A���V<7���\Ĭ �����W�m(���OD��' ^������D���@qy�T���1��Vo��X�+=�G"��^3kg?���<�r	5	wO������N�z������KX��B���ؿ� �KG�/�tt,\����wO��{�~�����p��GB�h"@Ae��E������Ə>d�5ƶ��x`��:a��Cqo=V}�:���b��W��n��X2Ҿs��x��ѣWOh�rՏ��4��B/�Ìk�X�p!v8wO�S���୆�_zS&>��G�����^#��[�%���m��q����U2��p�lW��liٴ]�pj�N�
��2Bz�S���Q��aeW`��᷿����XP��a� ��q�ģ�>���	a����!�l���F�f�B��q�u�4�$R(�6(�����e0�������Ъu������U'W�1�*�@b;h ��G����[F�ő�^�Px���j-��x��G"��.>�z^��L[+�f�&���r��FM����^���g��]+�懯�	R��*�m���ǟG���#��R��8�X�r%z����M'\����Q*�D�xyc�=�|�8�8��;�A,=�T���j�AJ�	P�N����0=jpu,0�L{�ء����H��fx��<�Za/DÇW.��ϡ�����FQhCJˢ�q��S��:)GC>O��j�	�x��'0a���ڥ'�H ���͵��@{.��+W��_��]�r��N�8�l3庐�}�I{8���Q��1�[���U�db�*h�B�3�-*G�1�߄��,����,0HhA�=~��Q����S��tX����CY��y�V$�~�N8nW;�(���P%aHc���3q��Qߩ�D|�t�@L)_D"V/��_-���O�F�w�L;H.��6Z�"�l����n�8�0�Bہ%��}�H��|Z��f0����m��OP���y-?��~��D�n��$v�bl���X>���]�{o���&��ke��ʛ���?^�xʑ����#�+#��(��T��r��`���8�����s��%?@��{�K�>�8����5B�jS���QW���1���a�؏'�߱��=�=v̙#�=��(Q��{�Rr�)W�����ĳ*$�:(�tۑ^�!�~����}��-$�$f�������Zt�^��rG�������跣�a�FOk�҅M8o�i8��(��$F\5�8�~����6<�23���ZEE``���u�l�`>�;c�8�h�P�\�IA`�!R�
}]
t8�!SJ����k��_��d�r9�{W|��,\~����E}������NҶc�U��k���w�{��B���I�
� �+�b����8���p��g`]&��:����{�r,�2�vĲd,`�HuY�%��m��]��� ��A�;Օ�S`N�V\��22�Pη�q]��6-��~�4���#q���ѥ�u��#T%Y5�<�����ѩ7.9
󾚋;@�/H+L%�l:�5+��1c��1�'~]�9�H%��RH:5���h�
泂���w	�=*>�e��g�
J��t%�(a`�e��u6�'i�C�
i���
��кA)��d'����2������Q@���I��!��a��F�iL{�>���&��=࢑���/�`��v�C�PSǒ���u�n?<Zjg�M�����������V�0�-��7^|���S�}��]��N��9}�Y�2���n��V�;�'X�Q*`��X��X�L$�<J�s���;�`=�î���Ʀh-��࣏��Gg�b1�Z2�IT�m��W'au�Zlק�N6��Wd��G�.G��.��d�D	1xAA)�TT���d&"
;¹�-0��v�bJFd��� ќ��G`�f�+ۈ;&� �}V�{������4����+��@�����|Q�3J���I����,D�.�L{�k�d/��o�E�a��M��(+oڍ\0����C�S.����Y�F��\!)�%EAS�#�+m�����(���ˮ�QhDz�B俞+,> �g܃~�C!�G�U�l[;�S4��3����1삑X�p`uj��ǀ��%�h�+��U���f�N�� �[�wQ�����dE8j�P���Z�m!0�T,v�k_�Ppې).B�!Z�Y[�̪�X�����y眂�T́S�P.`;:��툧��vsXٴ�~_�nB�� x8�2y��6���n��B���6�]��١��������1Ó��2n��u*�l�9�SB*GG�U|n�+��E�L�$	�U�as�ihI�E[q9KC�n;A+���䱦1�� \C^�0{����llhX�҂�\y�qe���>���]Q�Q�Kؐ��"i��.]�"�̒XT(�f����&��VsW+�Q�v<0�+��+��E[��h:ׂl�
;�e��)Z�#,� �~|/-���6�X�0ӪtA�����F�^�D����Э��ր����iȕ��PLCגH�I��d��|^��
G��#c���Z����
�o���f�^�����@;j{ht.2�۾ȱ�c¥�L�J��mH��D��Z��8VI<泅"z��߷�[6
���7ÉU!����T���D6���DcLi&�"_-v'�B`�9�#RKӨ|�K���۽=b�+�v�7�9���T���*�"U���
�S��x"���FÅM�����~j��6�AP2���O�B�?yM�v?�Z�Aw �MP���3��110Zڰ�?�*�Q)�"��)4/5�Q)�b#�klx����;���v�hȣ{��0�N(�<z���s}t��Kp§VƲ��E��o��Q(�g�$Cp�B������9�)�U_���}�U��\}��8tQ)bP{ID��D����E# �t�b/4iV�I�����X��Ac56l�H?e�U_�����A�9ƛ���Խ�����o�D*4�����pp��;>[�s���ɬd��=�|��aL������Z'�F
��gغ�Q|��@�$p��t@�Z������lJ{�$�o�`P�l��P�l��'�B/:&��2-2��kCiᣳD[AFGb��o9`E��=����M]T��),��;u���g_���>�=EjbP���o��j-�w��0�[r�9�L�Q],#J��-����!����4GQ ���b	��B�RSW+�B8g�l�Z��ܹ3L3%FB�%~��i�02)�LR(%�wa۴ќ/���R2��:\TY6�n1��(}��%���kW�8�8���o�Ըtᴣ�H2���>y��e؈��2�I���O���~�[Q�4O��	q�h�)�+ތ�C�,������$�P�QsT�D$�P\\�pMPuȐV���S�9�����C5/�s�-�'R9��I��0ۨ553v3bR뛰z�cF,�{��vJ�7�XDb%������5���u"�I3T�E-ơ�_q�B٘���Js�ZE����AnڼA���:����P��#�!)�lK�hD
���ɩ�}!Zr    IDATj"��ޅak(� ���ס�<�v����F�c/!����7p��kP�ұr�؆�g�G�ye�<|�2��4B=�<������'� ��,4r���ي�Fi�JH��b��%>Q�{�LD��\C{��Nhs��n��NQ��X�r�[��1�\V�%���ka�E�b�'�iH�%��d9�>Ǎ^�sRB.���dV�#4��x�韢����	��nC�bT����Cc;�,�:c2�XS+!0QR��c���Ii�567H~��f�/"b���J�4j�E}�!2T����F�q��Q	A�sX�z��'��ٹ�lh��Z��nM?�yZ�?�������n���x����\0���#.|��y�`�d~��76i�1<T?ŧ�����X��3�C�V\,�Z�J�J֜�[�3W`Ř{� H�UIO*��Q�$HH��,A�����4ũe���:�*�'�YʑV���,v�s���p�5ȥ�F�q�/�7��I�T�7�ݧI�ք�π���0���Ȕ�"� �7�2!������	�u�X�3YqJl��V����6��L���s���Qc��7�q�K�2�48�V�4n��:���S�d�l}g4�}	��~�.�]:����?jX>��^z����{9�ҩ~;x�
1.�v�6c��?��g)Z�L�l;����u"���w����X��I�.Z,L�b�Bj�^��d&I�`�F�4a����Z����\1���Dah�G����D�����%�6�>�c��3М��J��[�y��4s�&��_�Za�%D��8��r�bK��bPI�Ee�C]���X�'?�&�y?�kN8@���0	��g��(|�7����'����"�����~=�{`%:����7�v�[8�2
5c�	�o��g�P<��M�بu����h�[x���h��v���J?���PY�#q	��Ɯ�%E�J�j�>:�.�.c/@"!�R��"��1�o�y�B�R��\/'�=���>�y���͘N�3����<�*lF���N���n�ZcU�2�A߃�*��GEf�al�S��]�*�`1A�B�)wV��$���/f࣠�R<j�J�ÒԆ�S��N���b��	�ϛ��	Җ
U|[�m��`������q��}kW����@mFów�m�a,}������Ѝ2RQ��#���PD�[? 6��C���,d�<����%��5��kV�԰��.�?��E�+�NW�X,�6-4=|��&T�7�ȁN��G�c�^]PW�UR��:	]�g�a�+o �Wo�U]�IYBF������Z%�#�Ym����kk��� ��л�~'��f���	�p8 υ�j���EMW��|T�5_��";�:�ݫ�nb���@�$��*���B���$��T�(8� �9���C�ք�����3�ǡ�:I��n��,�nC���}�p��*�}�uq�lT�����x֞=Ʋ?�FOX���/_&��je�Z	�pa��3"�׿�w���͞�Դ$l%��i��E�dS#���f���S���5����a�U��0(�+�S�j�ç[��>uN�t5�tG�yr�T,Zp�w��iQZ�q]rz�6�N���}6����񻅓1�4�ثtS����*\�pp�sp�)g��r��.؊p���a�O��6��w��
[����S�#�D�DAY����P-V|�(?��
 ��nI>U(�5p�����bOĤ&,�P�0$f4�]e�%+_�߆N�Vl�`%��9�׌������6WF*��>��^_�A��$�}�s\������|��vH>������4��G_~���
^	Y;�XD3D�����_nŃ�_�BQ1�f,�b���m.��q3N�trF-�������Λ-(���g����?ؐ���ޅ�_~���T���E�1o�$t�I#�Pq�D�lW����&_�#�}>r]C�����K0�dt�Tˡ��&�ob��M���N85}��Mn�Q%��|"�闔G0,9���(�K|���1ĵK�h�Q0e���p���H�n�H�͗C�*dZBHk�XT�_W�=t�Aa�:h��H�p��Ǣs]=r�2�ٯP�:�G��g�J|��5�q2v��n۰t�{6��~��.7�_w�FI�D�M3��<�a�5���g���y�����Y[��r�J�̽�;�Z4uȯ���~�hDl�H#)%Ib���ֺm��{pԴ�تף�^ċ7]��7�E����x�#]�@Oa��Y�u�w��_J�X}�E�oҵ[g��s���=�U�Kf-�~������{Ҍ��+��bpfE&q�
���5O��-[��E�D'����+Sb�J�a�e��l]���b|�{�y�'2Vb���f��H ��BQ�yL����	6��'�|ad`�����ա���oF������8h�I�_����ƍ�8��Eبգ�
�vP�-�P�|��>�w�0�Q+ՉC�t���j����믽�\v��m��-�_�1n�5J�V6l�#�"����<���n3mևu�E3^�w���.���$&�R�t���ԫ�����A���Î�xc�EXx�t��M�C]��G"�9��%8�ĳ��<
[�l�c��Z�J}��N�#<�[֭E�#� ��3��Vj��<��	�+��V��Vd�w�w�{�%C���B�t��;�e=�7�c6M�m�nwjPpT�>y���M^$t�/�~y��ym�J����GO���._��Z�f&Fa�=�ϡ�����"}�X�a�)��]T(��[p���PHw�֏V#������	pY:<^)�k60c�8|�4��BU،Wg_��s�a�n�%���d?�UDhW�҉W���磴�I�Z^�sn�=�;�*��I��N-.�6O=ѾG�!L�$�I�Q
)��X� nhH.�a�Q�t-:�_���q��:��FIr�\�l���Y�ɍ�E!��0!���L�72r�U\�-�e�����'� �����+(~�	����v���>��1q�Ͽ>n	���a����&�{mڀ��e|��p��W��K��b��YC�N�'N���hX�.�=s��8yW��-#�P�t�R;e.6k�P�f�2�GX|�4�����R�F=8n��3.�<�>���Kxe�0,�?��v�N�&�އ ]���N<��ǠĘ��(Q3�J�LA�(Sn�LW�����~��ʭ��3ɮ4R�@�XϬu\�C��r��%��]�N��Ft��sa���"%)*�3�JDۃ�?;�,�>��g�dt����m��.nC����'~8z��=�ipI�5�Z*4�4���M|�?����Q*�15���i���<��'8a�Ll�jѼ�cl�ۃ�9f(���S����G���|ڈ{ߏc'^�u��m��6�_�����W���^���0�;������(d5/�5WL��{�iS�̇�a�Rȕ"\y�:��{�-A5"�J4\y���K�xv˚�Z��m�6��P��˔�Th,,ɧ.#�$)��)ZN2"߳��+��
nYVa:*��4��_�(xe2��]jhȗ����ݭ����t|�<�]<v�e��l��۱a����c�;o�h5v'5A�YB�¯���3u�ƈ�(T�5o����/l>`nLшJ��{�V5fp������BԼ	o, h�8���
�2`UZ=z����m�[�_��f.����ZD����W�=c:|�l�PҪ����3t�غ8�Bd�
Bt*7��\4Y�$�F`š$�J4�����.��G� jvg�3�f�r'K��L��<�"�4;+�)n��?�5<RY[��v7����5,]0��=NW���������Ġ	J�^&8�q(��P���?����,� �˴�NJ $,�z
�Z�����Z^�]#5|F/������k��B��b��.e���]�^N~����2uxF
MZ�T-�ЭC嵫�5}��r�8t����G&�$qR03u��Z(�5p� �\�ݨ��ƘGY	X�|BW��=�X�rv(�L&����Z��bq���L
㲶����cIӦăI����a,�n���Jsg5��R�� mZ������%N�a���m�7������?z֥��=>x�]j�J�P)V+ ��z�$��5$Q�y�� ����N6ZaR����
�/!��?�S�%�)Z��$�/�B��n�(�l=]*
��tRI]G�L�͗$�Ϧ�'w{��1E,C,Sig�Q�Z>|*7�z��H�$ϰ�h�[BZg>	P�N�B��������\�<ߚ�;�bi�x��}$������?��vJ������l�ǃ5zv�2��)�ѫ��)��B�h3�q[�1��ѳFL�����!1�x���u�,Q�T:��H���2�ZYk0����"�mnCJ�0*+v|��\��i��Ȯg I$���d��'�?G�ȫ�	��l�0�x
(D�{.��O�0� 6o���J>�˼Df3>0���h���|�L����K��tV�	D4��PG�v�4ĄuM[��wx�7�F	�
��l�K>���x��sQSi6�dh�Y脍b+�_1dԨ����;�Y�c�d�Q�[�j��6����6�%�i2I���>X���y�]J[�P���q:L�Z����BX)n)�n�˓��SKOk���؅GZ-�/c|�|/�&O�f������\ض	�+��<���m�ek�^��h������j���吧�x�>ue��}ʿ4]YT	�21�c���'^��_٭a�}�#g��<���x�3���5�a��C0c�.��.<�n����)W@d�ҭ�}urwuch�,�q�Γ��U�R�N����=Rv_=q�K�X�R�`,'�a��
����t�e��'�g�Zm|@��fg	� =m��c4���z7�C�b��7%���6e��R0p�$��SQX�+r�R˴�|^�x��7_q☑C_ޭa����3FM���6F���-jq����<{VTF�U���&|�H*a~�'�8�e,�[&�q,��-����8F�!-��	W�Q#���"��ƀ��7QCU��)i�/�I�
x�~�s:�*oD�zH���?�c�����<��3�ﬅNT�����P��7[�<hV�
Me�����Z\��E�b����|6/[8�ї���=�#?5e�/�j�"�a�mM��r�FP�4�ӷ�C�k@�cI^ �c�ſ��������?���RS��h�x$�Lx�\ghе3IV�Q�;D�h1&bw`�=�1M=8���֎���o�m��""����@I�3'#��.�� ���vu�c1<��lGr�b� ��ѱ��p�K���!{3�2�7�+	��BI�1b��-[8��=�RQ������d_�Ca�f?����x��@����m�k�3�J�.����s *��{��VW���{�L�N	������x_>V��P֫��G��ʆeo����R񝯖������\8Z�oy����,r0�&�RA�mNUʛ	��cP��=����8�(J%��f5M1�7W���Ο{��R	1�1�'Ti�&��r8b��Cy�����,���*!P�,F�W@my^�c-�=��0�+��R�mj،��M�&O^e���a5�C��5S�'�T�?�\d�U(�K0���،�/���D)�/�����|�7^!�iIN�XLOb���n X{�� �I �A/lDgm+�����=������ҵ��0�/b�[����,�vVD�c����������{$��'ޗ�O�>Co��ϡ0m��C'�u�-�j���0���%m���w[C؆#WV��8�d�E�]dc՝�p���ثc��^� L�����T�|�t���2�F��'(c�c�<b��8z�5�g����!й�A�+&�1��b	l��3)W�򐽗�߈��F<s�L���Km���`��X����`R,�*���롇��F���;>r:�:�ރ�/�OY���%�jh1��;X�%��b���F������=��Q��������0BW��$�e�ni�q�=w"�u�W#h�{7P\>b�T4��Wk�P�� �7�6u���:�z!o�IBC҈S��\5��H|�Y�Ӵ�����0d�	�]���ų0n��8f`/^I��P�X8w>V����D�����a�3X�a�~ElT�qg�!L�@�h^�}\~��i'��0*�mhp�f[ҍ�i���7���5����a��I�֩C�W�E%��KF�P�9�N�����u���p264E�b��8b̵�W퍂Q�*$��\��R�������q��&���M!�`v�C�h3�_2cƟ�c�F�g#O���ebѼ�X��[r�bt����܇|DF�N 5���GLG�����`i���=��%܄�w��0dEqʜ'��1�&�0D��E���T�(,�3];w��^K��p���O��N���=dȉ�B	�����3�.�c���Y�����z�l�1�I�]�<ŗ5A���v�n����DegK(�d7�&�ml����7b�*���T��[��v��y�Gv%����2��l��X��s���1i���dInO���<�J����U���ѹs�j���	�K1BF{^C�R�95e��,��]�|�^(Y�`�Q��	A`�K*1-���~��8W%���zzVP����%31n�98f`_�0�"<±M,�{V�Z�89��'�{�=��c؈��}����,�P2
s���u�s(I<F�c�}}k���h�a��C	�1�4��蓙kT>���Fa�܉�Թ{�����/�a�㹫��x���t��]�u��rfM^��hJ��	�gF�d��c:"����� {Z��C�a�2�����lØ0�,;��pl�*��[�Pr�\�JA[ƞ��#>$a���
�_(�q=�8�������+���y���2rҼ?��0T��鞮sa9�,K)"������F`��ɨ��M<���ɰ)�#GUB	�4�{����O��KGHKPTL>s�O^�c/��l/�*��M�����KbY	��'&�_�0,;�\-;(���9�_<��� ��%M)��0eo���j�W�{��|.��JP��a#����ֆa��v{�6Ɗ�;y���j�a�a�^=�1T��:�1�\��2̝;]:u�K�{��#b�h�+WUɨxs��Æf�'-��/��L/A��&��$S@B$�e�QC��;��v�-ư��w� H�)2�j�~�B��w��/����$��m,�V�z'|U�=��r5f
����/��.إa�Y��QUI�p3V�qyn���C�8D��G�9b�ܧ�b��P���Y$WFd6�mF��1��l:�q:�Lnd���0��F��tT<���Y'�de�7��s�i8��d�@� �|��}L��z�8��ӽШU#G!�te�k�#LH�T�S�J8�a�T6���vu}��q'�9���L&��،��zl�3fa��q��_���EQ9�O�馛��悔ޝR(����~�1�8�7l�5t�$t?�:�z&FW*��8�!��k���RU$��p�%��vø���O9yޟ�j:�N@.��%�!�/n��gxeŵ����9EN�"L8p�Uh�7�?<�1Zݡ�^E�E�
A�AK�n��à��(,���	��&V��o8�G���(�(h\Z,�{5z�$�P���k��P�ʎ��ŋ)#QH+5ZQ�$��8�r#:�#8�6�����e@o�ۧ^PhZ��]�^�����o���JV~�μ&O�����=G �+W(��?��ngM��� ��p]�7$���{�kk�1�m���؉�L�����$� �M�8V��	�x��o��A�l����2'�B(�Co}:c�
�o�M��\����gJ��􀓿-]��⺃	�
ƺj�1QT����I�P#���![�c���H`}
�����l՛aI �Qqh�z�    IDAT���_��@�d�-\�����m~�GT���.D�Yu�Bz[��T[ �:�u��0k���|$�&���0�$�4/_4��=��v���q@�d�+`��}#ȣC*@��`��HBƜ���t��bHJevo�sۊM���Bj��mo���Dx�03Uȗ�l��I�0��I�������A'���+��Z��L�� /@п��U�CgF���/�1#�V�^!}�+P��x�3�*q�2�
~��c�^��A��Q$a��g	L��6�hv&n��}XE+�Ð�Wo"M�,�f���<�F"x��͟�,�ui�E)��ga!�D���#��,7�\��!�/�LjP�CGI))<]�O!?�0��&1 ������)gU���9�{镴r+���*A�:4M�\�҈i�g�[H�j�c|��j�ؾ��g�,����6?=!#W��Ie�FI<I��\i�q�;k�|��}��F�rAC�)� Nt�Q#Ur,ͤ��y��l��(��%7���![�fkP���?K�6�} �t�pG���2'�݌�܎������??	I�)����"�|aK�Q��G�c;!�8A�DȈ6;�b�x���R�>����+8"��{��q+v����x�$4
�z�X��uJm�6@������0ڄ�jWUR1{Ob�Z�Qw��{&�+�2d�c��I���Q.Tx���(V�� ?R	�Z�yTF�����.�X�����_p����l|4��7�#Ij�O;i�I�T1�ib�\�?5*{�X��%����0	K���(r΂iā��(�[b;3�؃%�n4.A��Z��\v�lE�m0�ۨ0���+�xbl�c(�yk��&�h_�+nq��i��#n)#����f�Ҫ%��!��̡x�=�:�L�S����Gy �V�^*���X̋k%��l�k�ZO��c=*wGMg����Crbe�!�8�I�+�Y�0i�'����sɼDȢ��Ğ�>1lz	~�xO��U��k�O�?!k���%��Da ^)`4y��z��%$w��hLP�x����7Oo�-q��J�t�+Hnl�	�I����O�ѿH-�<�J�8�����[��s���-�S~�1���l9^Ib���mx���-�ɱXFȄQ���v9ȚG쩨%ƽ?R�
���q�{'�xw�bj�4}al��"U����h|��]�֯����cH����ю骂ޫ�͆��bɆ$�'#n�8����$i����\kI�*�H������_�Ժ�3$V�5�0�¸�&�^�k8DV��	h4�c�v%�xr���Q8��p�̟a�+y�R��^J����7Y�ja:n�����!���M����r��GM�G|�$�k���oF{��u�j��Ee�-E� �zc���B0�`�Eۑ}ng�۟���M$y�� �a�?B���a�aҕ���G��� �Cl��&qd퉇��J��1q��i��ai�����~\�R�Dr8Z_�T9�G%{}�o��j �S���{�>Lؾ%�r��x�v ��tQ����j�I=%� C69 |H���sw������#_�8f2]�ױBH�[�Z�&�=.��	��!���7��"Yud���?�*�/���]hh�5�RQ8�T*\1�������D�5)��sԿT�Ί-��Q��ѹ�����i���%� Kj�4��%=^DR��� �Klb:�|���x�<I�J�h�{��H�2C��[��S1h��e�P��k@]M��7�(l�WjĖmM��J�lMg�k:	�g!�����0"�?[]]YH�]=$Uٴb⑊C}�@�Z!�X�������
ٶ}v����[�ў����D�/u3x
�z��E���!���FO�|�r��b-yF[�dL/�=���Q���lpe�r��|Ԛ6�}�W>|���V:=�b���PW��|�lY��"��s �p:����EIKAKנ�(p�>�5�@k�QM҇V}�=>�V_�ŃQ����`_��a���}G���2��˜C@0��|+�B�$S��M0��	>���J�RNO뤬-��g�B�LF#iH��뜩�ѻS5>~�oX� o�N�C�9��?2�(����T��o���<�L�|*`T��w�G�����ed����2wQ��˅�(UM���V���*��dUA	ͨ܄��%�b�P@�<�����ٴ��5�$g��)�+w�U����ln�)UwT>/G��IC�|�q���m�z
��ADb��ql�?��*-,�n8�����r�=��A/�?������Ko��OEV��hI`��#n�y�o��\���y	g�v.��0q��[���g`ejĚ*�q�h��jy�Ʉ6A�WtYHRO]��=(
�?�+Ir��*+I�e�̕�Lg�/���wa)�9�P�V���/.��'P���z�s�L�, �ƢIĮ���� r|R�U���^�f�\�V�JbFd�7�ؖN0INI*�5�%��n	�TVi#��>���/�A�{��A�^��|�����8J*���x�u��w�Mx��_��3�g�ES�F٠�ԅz�Xצ��LZh��*7��L̻U���DtԷ�[��͊m�u� s��?�.S�(f ������Yp�(e�~��$6%gUj��G�l��앴u���7Q��B�D����	�1�����q�_�~{w�
#Ij �8VUa�B|�������Kg!_u0rf�����_�� w�L�M9!ZT�_:��D���t�6���3p�����?�S@A�n
��KQ�����c��]�#�&��Il�\ ���ab������p�����썜Ü�BT,�4�� i���B"q&$ơ2 �2��HS��o~���z��z1��W�荰�֌4��`�y����t���+f.�~ρֽ?"�k�1H�Cq������q�=YjnSK�=9F�㎉X2
:v�(�x�iȌ�;���ΤMB��0k�|{��(��-A*��ܹaȅ�E<�� �����b���~�c�d�_.��tQ�	��U|�e�Ðe|�ylj`�S ��H�	�-Ǐ��)�6��}�L�N�)���mt��*aAP��(��sE�.�QS��m�]3V��!Io��~G+,�y��T-�����a�x����w�1Sh����v���6�q���׈I�~�6�N�<�mKf�W�[#5�	���J薘`q&@��isp�%W��?Mz�"\߅ǐ��������۫�����_݃O��A�=�8,�,�>R�'�$7R{a��#�SÓ�2��m�p��9_�*{�t.���vE�PVd�%�?(+��D4QRV���e;C�� j^��<��*��x!�8pX~$�y�XK�Ca�:���F��}4W<Fblʩ�u`��6������NB�q9	�j9s��@o��L-�{
���l�b��K���>�2Y�yD����qV�9���c8���Qs�D��hLt�<aq���0�fv�K�{%1U(O������б8�F�kz��;�H�J�TX�e)Q)x�,qE�<�����̒i�l�0֯�0�����.���Tʉ
�����𑳰߰���u���a���ѦPr�̾n��o?�I��� U�lI,�t���\u�m8���1�r��̮B	2��rR6B7��Q�������{�ۯ/�(�u\��\�����4�*M6��(�"Xr��u��1@fç܀��y�8l���,n�U��T�Y�HJ,)�w�Ie��ft
?�P2��0�O��&��S���)�:m[�����=�&�z�TӐ�_B �r�Ģ��S�Ю�+7�[�ᔓ���C����7Pg����&+_x���	��`l�2�T��0X	��rK�2<8����W���'7@��,�=ߓ0��_@�i��f�3[��q�R�_�#���z���[ߌ��"��Z��\K��e�Qs�Ua��a$ɧ��Y6P���Uۀ�,��C�; ]�j,E�O�!S]+B����1��_��E���F1Jn����F���Sy�Sǎ� �5-�(���i��
��f�N9Jw�c����CGLG�n����W%1�"˴z� �ӗ����!,}("�"qMv?�u��P�Jܔ�&Y�.RQE [�Im�F.q�X����<#�����G��'�1�J�T�'�妆p�;�p�1����UF\�)Ɩ7��7b��a���0�PE�43�|��!o�*��e4�������a�=PH�:@�!�_���ʫ�[�y��)�^[^v����&iZ��%�T��(Wc�3;�Aя�1چ�K�`@]�~��iP`�/5�Pq]�S�'��G�N����W�Jꪥ靌��G���[~���?���3�e���mT������d+�&&9Cd�&����ܭ�����!����o������,2��`��iZ	f���9Wi��%9��~��_�EU�e�%mB��}��?9i�Ͽªą�N����j�ap4E"�,t��`�/�䳇�ic+({�M���b�Hش8�-���dd�IL�֪z\T�4��o��������a�ᆊ[���2�ފ"�H�iőE�7	��7�9�R��V�4�?j�a�kS����14H�[p}�:d�?�'?�+������:eɾ�<IO�j�f���_�lF,�IB��k$i\k��˯��y�>�n|�Պx�n�BtO��+ K����&�G�v�fcG����X��4[�ߘ=���\�����E�2np%-��z���rو�^m}nw���� ��Ð:ݴ��`�l��>O,�	�;���I
�x��vx�U٨"_M��yղt˸[��Tǵ2���~��50�3�^�Ԑ"�Ꮠ@6�uGu8��jng��Ƕ�"Z��a��0�bzU�#+�j�P�/iKc��+��#3���=r���s�
C���l˫�D+�|H1�[�����n���Gc���W9��1�V=�u�\W�h�]��n
��P�\��X��/}�����C���Iw�!�C؄�%/��NƆ�ȑ�Q����+���!�ǿ��[����a4-[8��ї\��<�#珘4����0��Z�.�d�2����F��a������.?�/=Oe�0 �yp�G��8�`I��ۣW�mC��r�/n�Wf+��x
�?gMX��A��+�r���sD�p�:�Q&�9CSp�v��4�� �M#w����WV��/��6z���7O�Ƙ��ڭa�}����<�_�aD�ZG��-�v�����f6��o���ϱ�+`�]�d�Z&�n<�2)�^��*Q�&NB���H]���O��VǼ�Kqǯ^�ާO�'�j����/_����<M�`�(i��cH�о䳨A{0fh���?k�>z��)s~�V��4X���p^)�
�9E�����1�����ֽ{�Mm��}MҢnG��&Q�t��X
l�� ƥa8�٩m�H��6����Ŧ��Dyh��R�D=t[2���QU�s[r�{�8U�+��@��媅����A��4����C�Ƚ��%�S�*Q�A����
�����'x��Yx����l{�9=&�� �l��{k���Dmߣd���웴�iKF��n5lT�w�s(���헷�c����ᣦ̽�m�����M6V��i�BP�����;�G������o��x$wi$��ÃκL��>e���,9�⍕�t�yʓ�G���-˔�J+�����r5~�ԣ�α��� K�jx&s3�+Q	�a�Vj�$��S���;��:<Ɋ�����}�ހ��	������ݐ��M�jn���H��՚QW��,����z'5Pn�TO\�;J4��ka��n֜}���5U�W�}�7�]8]eK\�z���a�(�勧}�ҋ/X��P���#'Ϲ�-�����DÐ-3f|&4K�Ϸ��Ƨk^�|�����X��r��ϛ�a�Ð�;��Q�Tqf	�o� ���v�� Ҝ��O�W��7?^�,��5ٕ����H�u��Đ��7������rr{&I�QW/�}\���s���Ƀ$S���-�TrT���
!��(7�R�6t�>�SKf⅗�/��Z�Y��0"2*aek��{��Y3Q���C�J�b��!�S1S������\y����ڔc��0����`�.�*ӸBHè-|�ՋG���b٪�z�soCS�Y�q�z���o�3�^,au��Qml�y��t�Xh{����T,9Q��]�J���t²ZLՠ�i+:�BT����f�/�_�G�2KpP�c�	���G�1z����W	�����Z���ۊ~}���.�N��2��9��ٚ� �S�D�V�!�C3`�[ѱ�!^�g6�!��5a�|�x+np��#�$�d_�P���OB�3f���a���V���=ޤ(�O�Z��T���e"DI'B]�#��e�؈����B�Th�a���������/���� l
�����ceR�Ls�!��-"]���et��	����Q~�Y������j��: 5CH>Bq�
dGa˓W�*�/D�� �H�N�JRړ�=����3�l	2��!j�D��8�op��*�@���FM��ن?�t9�"˸(�}|��L
�|c�Ks���g�B�ϑ�.׸-�V&x��R�hO���,���2s�'+/����:�Z<�&����K��,)S��GU��l��Tl��<�F~��#�ڧd.�1NL���������SK�3���F���c8吽���"<Q�Z��
����Pf!RnqoCT�X��/gl'{ �����w����q�������1&�b(~�,��Pq~{sk
gz>JhTkE�4���V\�	��1��E� ꔃP#q��b���Y��9��Q�x��Ͽ�^�Ǥ�VL�~�b�I�<�%�����^à��*�(q���,���닆a�3q�atw6��Z&.�[�a)/�O�Ic�W_��OE��`4���g�aPK��t��R���Mq�|3�j��{y����?�+w/�/<�/���g>{�Vӱ$�y���J
 j���Kzs�҇0�y8f�upS]QD5�	�m	�!ق�y��D����Q�����fb���qD��Đ�+���(K�Ͳ8�[:硗LG���
�g  XՈ���0V��M��6b�ڒ|��ÈҒ ꑇN�:���"\5c����2�l8i�\�@ΦӢqFؘ�0sҍ8l��(���?%�Z��� �� S-g�<�n�kR+,*��N	G��1���Y��[��G���	�(R*�H�cW[����\5����W�u`ظk���?ǠS`v�m��HO�H|��4�H�����������:� Kⅻ����g��=��q�� _R6:�Ӗ
9X)�G�Dߋo��c |�D0�����	o�R��*�l�a�ݎ>���TʄdV4hiA*Q��s�+]�i���!��E��B l8���{�42Ӭ����+P�P�b>c�Sº��wPnB~u[})�z&�&��CD�Y�&X����ۯ��?�í+c���@$��ċ(�:�PP���~Ç�:��#�Uݱ>�ê� b}��x�����"nC�e��<^h80�[�����2�ǜ�c�)�O��f�N5B.NŬB4,'e���	�N���X�kx�����H��ٽa�Rs�]f���!Z�:��8�'U��y#q�vXF'�_<
�ǝ���<����OJfˠ�L!W��W56t�C�,�����[���V�|4�q�3�D&�Ze�N�@JREt�����+����2#'\��:�uA�\[��:��/���}�u\q�B`�����#N��&_�Nu�rQ���0����h��C�dJ������e�L��1p?�,�Ejy?R���pH�����G�B��C�1PV�Rg�$�D�uC�-I��-����&�Xq�CGM��`[BI��j�ֆ�	ʨ�c��1�t��8f� ��BK�p��zI���L����s�V�~��<|��}���ʴl�'$�����Q��/���c��*��	��6`�'�b���QX������_��i+���y�>�Px8�>��C���5hU��T�@L�    IDATv��/j[�|YÐ�'ӗR�ݍx�q���#���n�t��?�I�R�%�w���Y���л��KY5v�cm�|2�n��ضy�{�o�-�6@e��j��*܌�n�p�@�Iy5�F��җ�q�&���b�������y�NZ����M�v�N���d�@�i1ތ�����(5"��r���I+�a�6��W*ɺa�_
������ �,�"85]��)4�
"����YxLwiINQ�!�6�e��uQ���f���f��yU��'���
b��oy�3�j��+<�I�#�DS�uh�-ø����9y��m�I#�$�$�gV�#P��6j-]䤂����#���k:�.қ����0�ڽ��7kD��8M���1��*E�|~���.I�uN�q5���eW���Dl*�(-�2[�wcU�2�l;KXI�H�6f*��\�L鴃b!�T�VDg�b�Ȏ4K�)x�D�7 y�������G��v^A���0SҊ�����Q���l����Ɗ͒����7���8a�x��?z�Isi�aHqse�9�/]I��V/�aK�wQv}�p�TZ��n�Uf��e����7��s)�M^�@�	U+\���0ĿDj��xϗ)-x�Z�a�@x�Iƚ�����2%"|#�J�*��jh*9qY�����%�({�+.SC(�)�B"��i������^]�2T�`"���҆�D_����0�4%�,J�}��P����/H��F������E��l���\*�o\�p�=�1����Dn`+* �x%�)���[�JV��(���I-#�c�z�W-%��7�+aS�J@��@�`�l�/��YJ\���c�8�Ed�iY�XM�1����lPF�hq]�G7
�!��s�َ��[P�'�<d3�_c��-��n�3��=��T]VAɲ��	˟���YK6��G(�x��j�RN��H��*�P��(��0V���٣��{�����"�3,)����Q��R�,d�Q�U�M+Q+Hq	�j�t�|p�4t�!�����K�-���*�)T�.%���ϝ<��|��z�ghJc]QI2�(�6��&�@,+��Mtۅ��W'7�"6a�)�*'o����s�PQ����w��~.{8�c�ՠt�(OxL���*I���>��-9���B��)U򲖮g�c��0��<��6 uڮ�|�����yLɖᯠ<]�Cn %���{�*�bY����IOD*'5�J����I�9�O���I
���~�����8�I�TU�A�'��.zn����JA��Ϲ���8�5uSI>p_�]NI�ZA�c2:E���U6��A��[11q'��/:|�ra��Y�}YT���vF	;�dُ�eΐ�0�ސLSe�[�S�>�T�J�/���=��ۃ.��$TJ�"P8Q-���"5�u2�(�p]��Д˫�C�k��#�
!��Qln�ϕ8 �R���U�r�I}c)���u't��l�5!���GVg�Z:V�_DZK����;#W�s�0*
קw��`%
�+wI�It�p�M��JjE'�	p�����P��KlYS�_��JO�PjY�đ!��,�[U�7׀�AI1Ű^P�l��Q��N#�z�����qJ���W|��A�("��bI�%���dm���TTjB�Y��aC`��pR5ꁺEX��M�$E������VXB�a�{�Fs���	���<)���q_Z��Q�b�,-M��*�JY�dYF^N��ٍ�A�.��r	�Cɍ&ľ��d�#>������_B�LŇC-.�������+�oǥ� ��j���-t���lM5�%5��$��D�v)�3�BP'�7cl+�<�n I�%�r�H��������D�c!�J�c��X� D���*�8��\��ݺ�Cڑ!N�4:o�/b��*E�y(�s�i*GH�����|^Z	ZA<�DV+N�K�	�S\��+�2]�d��=w�l��x^#,ǂg����&�i��\��|N
�b���t�A)�jH-V�|G�%a��'�����Z:h��fb(���$r6+��0@���s#hl����,XF���Q���"��(A�oy���k{��C��*}S��ɤ��,&�erZ;B���6C3#)b"�M9�BH�g�34�]��r*�R2m��!� ��u�䉬�,j���؉T@6A.�T��G(����t��ư#zL�y�"�� n䢙���� �T-rVHY)��y���#��p�ɕD����p�+8_ �+�'*[�Ԭ1|��,Sl'R<;L��������\��Y(�Bx�S�\�衐;��P,Y����0ڷp�2k�!koE���L`*3-�F�F9����7���	U�#d�.̭nIT!&#���pɱ)�<ܮʺi�2Bu�٢���"���	�R)�~lp	P,�^��Z�\>&�
q����p#���b�ơ�eSY���c��)4E1�t�B�P��R7�Ur��*�&هm[s�4�L#Dѣa8r8��Ӏjzٲ���PE"�#�@���K�BB}i�E�?�&���P�&�ؕ�X�p�W��P7 ���F������&��0��'aӨ��oF��	���i�:��YzU��CN�#t���e��\C���
��ѳX�M�Ig�d��r&2`���.�ha��e갵"
�m��nظU��u���T�[���5Ǉ����a�a���(����1�����Q<�L�Z���zҠl�% a�C�ə�B�sa��<�xՖ���|��W�P(QۡNr(�����\tѣ�^H�r��l]�X[_�2����پ���|*:B���b�Qx"��͓��B�ۄ���ǡ�Bm�Z�������+��ߗ��G(4n·���y��?�U.oP3��zϬ^O�@��p��4��طe�ې��r���W=�[��;��ף�Cg�|�x�w�A��M]R.z�쁗�[����c�늌��J���{���O�0�����*ui�������L�]Y���]�RN�����s͠���c��zⵕ���ǀ��q��A��^��	��� �WF��0��1x`?4or��k�fK[K��/ۣ�ve(��1M;i��h흮�
��*�4�f��_@��Ƀ:�_o�<�V�
|��s��n�� �Y�a�]t�i�k�:|��'0�4�[?��}7\�����!���%Nxc}�B�湗�i<�*�IT�KRjVa�bȡ}1qTo��%��Qk��o�����⋿���	=�6�TzX{�!�p�/q�Q�b�y=�֫e��� �����;؝��h0P�\��ȕ!"jϬ��pr������G3�E��
Qӧ9�����{�O1�GCq�`/�=Ė���l�r˳���p���!p��/oA���e���^�V"����Si�k�1�i��3NڳRs;�:I��ت�Oվ�����}�&e"�o�ms��+n~~�%�Aˮ=/<�1~���y�yx�X��x�ݷ�ǣ�OŲe/���`�Kw����7�?��&�u�,�Q�A�.�uK03���������O���4�P�fk��z�zv��o�}�æ='?�� �&���&�C���ptg�x����p�����b՛y���ߠ��P�!ym���zbA�"M덫���s0e΋�|�m�+��߽Z��F��� ��|�࡬G��s����Q_���?���A)@�J�>[�T�!�7c��Y�}�y�hm[;@Lڃ��a�a(JQ<>����5�,7c`�z\x� �h��t�B���ۀ)�5�t0k�Op弋���>��~�Щ�߼?�w��7�ޔHےK��-f��t�s�˿�՛�j$��������]0��>�A�k?l+z�ׄ*�N�����o��Go�����ƕW��{�1v�i�h�8��#q�{bܔ���v(P��C��o���������0�(����t���Ȕ�a��`d��Kđ}�a⸓1z�C8��� �ࣿz
MZ/�4�L��'��ϋ��{��#��R���Y�w����� U�EDε�+��b���G��`����� <����۶YI���Y�ڔJ�*�GCC�p�)��ē:�򫟄�aXv=����N�|����Y+p�Q��ck�v�68���#�����^�S�d4~��!X�6��~�
�N7ԊDX���Ȱ
�n�)͍ͮ�p�1�����p�#(:�6�[ؿ�<_�z�s8x�!��I��}�r�y�x���b��0tԷ1�ʟ�SO��'�b�5� �=K����8��#pѕ�0LQ8����4�SZAHIM�oވ>=:b¨��r�
�6T&���ߏ��Fc��?}���3�����em �~7�$̜r/>3{!��yW��,Æ�!#����c4ߵ`�ɗ���n=���>r��)s�i�a(�E����I����3~	��	��Maܘ�8��G����M�*�0컇�G�,��	L��,<�Л����ix�mx`��~��V��-�p�����5�g/�OwGFKJ2͊��`�-s��T��{�`�E=1}��0;tG��ѷC��c��ᓟD���q�=qͬп�>�1���ﮧp�ȓ1lگ��O��N��u7��:[7�ǹ������a3�v_�Q;�Twdc�8� ��G@=ִ-�qż�q�-´I�`�m�����̪�Z����93��PFA�!16�r��(j�I~#�Ad�� )6�WQA�A��$�2 خb	2���9gN��f�ooa�k�y<O���o�o���U�������ˮ�h�_��폂�C���hށUs/������� ,�#P�H"Ef�^R�j��|�;��,
=4�_'�|��lF5��&^��lĶ5�u�ނYS���;_⩗_�-�]���X���֡.�桤���؉��(�ɜ1���h㞧6�t�f��D�T�7�@�9b*sp߄JQ����s���*6�F$�Y�%[8nZ��8	���7O{��è���
\��Ӟƙ��E��;`���?�d465`�X���Wo�)d���Ty�H����$R�Ԝ<�&����8��/ ��|��qr�1�:|!�pg$lb!���fa�Ⱦ��ۘ��i4
:uA}���i����w�+Y5��T���dT&$;I�q��ۋ/����w�植�N��l��]9�3z�聑����{@m��~��x�=��e/B���j�6�\$����/C	���5@���WS�:�.+M�.��^��/���kZ�9�ǅ��":�U�:�L��7���=�`~'��v���D�;�9�~֯q]���C aǝl�R�c �,����&�M�g�'�OC�)1�@N�[��_����_�� ���8n�Gu������/�@���]w\�ʝ��-@^PCYɚ��G,�h[��A�h�b������?���x�<J��F�����>5�t&o7�P,��%e"VW�ӎ;'��S�s�lM��w߆�`j9��4qF��(������a��g~->(V
�W���슛H��P:�+�Ӊ��M=I�yU�����il7"!�\t�! Yc`��j|�����'�_|�vN�]���rQTt$_�ݏ��~�Aꯨ>���d{�
�
EE��A�� %>oBN���\��t����2�G�>��O?a�?I�L�`%�����X��Zl���d�p'��D��g$-��u[�O�.֌PN������V��c��C�0���=sU)Ȑ�=��a#�#��S7�7Z�P��H.o����Ò0R-h'�nG�D
��|dH�D�3
�$d��*�����,�]e���P�ށi���g"9~�$�k�!H��$� O�Y��h���:k2�0-)�x��.|2R��P��Ɍ�K�$�3$�C�ɢHc�g/�t$`D���#�!��`�a�`F"[63�8`��z:Ú(�t>Ӏ�hJ�hױ�Ob-[��Z\͖���,�WXۢ��j@E'������I,����S�1�%f�4$�..�O� KBʰ�H�Y��:dL��.)YZ������=A�I��_h����Q$�Is�n�M���1H���a�SU0�Լ�?�d�ivj�z���_VGtU�\�J8Sj�;
�J�+����룣��b�ϝ���$��}�D"P�xV�	^�t�NӤ_J�K�=�ᙓ.1��~��č��L�#E�J�%�_P\�I�E�uN�3`mr�9V��S��G �hD�~^i�����iK�(E\�J|�t��n=��A�Fe�!�q�Rw�J1D�#{�l�4���N��7��*�ihhDT5� �GR�<$�s�1�p�Ej��bP��$b!��4!�#��ޑ���Sy�&��V~��AR��X:}!�u/DP�{���1�5����o����͒2T��Fm!��4L�:�&�i@*�+t)H1UN	�)�����P;:'Ľ��� �cW4fd�dd.���E�r���
� ���A��X�6��,�6Gy"�VEgԃ�y�Ds-l"f�izNw(�����<�"��$�!��7�0�X���Cد ������)��Mք���@���}P5���BGSFB�{o4e迉��f|��+p��/�q�o���q@�X�xŐ!��~��u���<ڣ&b>K�M�r�B�I2����&Rk�L�KuDVO%qŁx�|�D���PvҁBH�KLx�� ���[f�F�IO h5��s�t����"<j6����oݠ
�C9��~�<xD�<��A����뽨�	(��P�l&Q�y=��z�A�
�����T>�z<*)�O�r��i� �
���#1�I�>��4�KV-wׂ���]�8��/�:�;_Bp>��f`��AX����hx���EZɛ�"�[�E��ۣ- a;�G���+��I�?�I�a,���&�@��rX|:�:7㍹� f=��`n$�H�o����Ť��Fd@m��Jq�)��QKF�ʢ-�w�s/n�!�(��D�R��jT���J���Sg<�rIz󎞡��AHw�^�g#�+�e��&�q?�W�+1֔��E�7�c2��G�n�@a�
}t�/q7L����B��F����z�|�r��@��:�o*���/�Y��v�/�NG��)���v�N��=Q:�UR�%oefP�Ϡ�ڃWg�dvv�}#�-qc9�<�n��K�N���'��[�#����x��;Pc�:͊
_��M/a�ߖ��i1��j���9�����<�j�1�aĔ#��d��1�Ɣ�]�{&_rݐ���1���l�]��j�=����G
���$��AnN�H"�I�����������V�G�hE�\(�&�i�Y�G��Q����
ӟ� w���Q��4m/e�\��#�nDAf'�?8�l����+�-"F➠6W���Px�(��	;��,(�R>z?ϣ��qB5bϣ��ֲ槫Q�z)T���\2��E�m�SN��~���Dq�	�OX�z���l/�^�Ѳ`��K�J��,��~脻l�a����]���*d��i�J�Sȓh��2v�0�ټW}�{@"#�%T���$��΁T����v3)�������8��(�[[!��2��jtqvc��I�̯�'Jw[���d�Fb2J)�.��ec��� ��c8v�M�����yXWI��9zқ����j�3��l�db�Q�~�M�DW���^�}&,D����L<�����y3'^:|蠊{�%+F�������`��#���?�\�d�t�eu�[
|��1����^5���9��AWE"o4�A�:�R�T\� }�Z7�=�nԨG0��x�i @d#���$�G�N9v3
t"Z���=q`� �m��N]q^RC��G���Ǣ�	�!-�p�U���*Hd��<B�6ȨLGF;�{�il_�?P�Z��G
�b���)
t+-T=�b6�|��a1���,���<y��g�gM�lXt�ڃ��c���y�bh�����2���
6��Q����C�l��b�s  �IDATFِͪL�9̫�O����nGn��ۓ,��	c���+� �H�=�N�)G I�*�]�(���3]�`q�a�|,-C3�_a��ɀ���d .}��%�qR��ИHs
H���=��-_����j'^6��)9����<N�x�]�tw�����齿b��_Q��4���i��B$'i��k�][��̀e�^��L-DѠv�ek<}�*���0��gM��"�砆�p��qC��5���Ὕ�C�C�TB^sg��BQ������nA��5�[u/?�{��*�s=��B�"���9���$ʮ��
���l}�ށ:�I9��*�àݤ�M��J�Ŵ����x�̀�`6{�7L�������$��h2&���;����|��)9���^,A�S����a����"D�8��]�]/-㬈��4HE5��KW�b[&��(�q�5�����7,F��6Iw1-D[�.?Ʒ�h�y3�\6|h�k���ax4C%Z1u�N��o.it�g Ό�ͯ�n�}�Y�����N3f݋�Y��F���rc3�=J:����W;!)繴��+ܹ P�u\�#�k�l��x�-�U��l�d�c&��/N�	���-U������/�~�0.����EF��`(٘���<��l1F.ZP��*�~���HN��^��=�P(���pn��FL�2ŕ�d J�:i�#�X2$��ګ�������ߑ���c<�h�ء����m��
�8�:/t��n�+��v`�Q��g��(<:T����.��nhsH'���Q7s f_�d��^툤�+��jyj͕�o����i �đkVc��[������N�8}N;����"5�n��TTn�r5MX����@���c�:�^AM̮�0���[B�(Ix�����a5p�̌�2p����ɇ����ݜ60��1"���.��	}&>�_� 4��<]�	��e�fN���磋W�:����b��9=e�m�l�@P���IL����"���M�~�Hv�p�6�{/��LI�SX�2"8��<u��q��Q鈔,x@|^̊~���M��l�#Ϩ��{ou=F���ɓ�3�N�͚�A�f�uL��fl۾�5�L�.���aPZ*�ἴA���D�{A���%a�?�]lM�㟞t��#77Eg���`��񮖊�j��c,A��H7@���U~ �.�X0{��MW�Y	Sr�H��/	������p����QQ0i h��a�z�(N����F����E^$��:{i�h���PF�낳�ގ�0Zȭ�}o*g*��pD~b�a4�Q��>2�� US1f�H�:�'�3ҀM�O�6_T��j!
.��ǟ���m��6E�Dɉ����.�,�� d�a���M��B�F����9�AD�~�-��il�1��[�j��`��`*]�{�c�����h�oo�2��0�g�E-p-\�l��3�5�Ԡ��y>x��H}�(��"���3j����>�OйK�)��2"]ݼ;V- �Q��������Da~G��I9��Dݣ��Z�;�N��af����
���^����yX'��݌\���a�vL�q��ĉpꩽВLs5����4m**+w����^� �/��O�+uk!��%�'�*hH��->Z�J1�~�<����0��н�C��8�&��Q݀&L� �|u���LZ�G	���[ܶT�@G��3'�f��A�������1d���:f1��B� �"[%4�jc�H)�$2v�8���EB��x�ILA�C��+��o+�[#���m��~��ܾ��& J�R!?JXr����Q� f��#�[�`��k`�<ͮ�1����(YM�:��D�8F7�pN<�R���ɓ��˯��Ћ!��oJP���#��ʫ�z�5�����a!�ɼ~��_���|���WCs��~����׎'ۉ�1na܈�P�[���,��g�{�Z$-���j*�-�د�x`L˼{n�p��?���hђ��f�;u�b�!�!���t�N.�D��# 9̚Gmwj_s���W��p4��+��ހʏ6��:���D�@e�4f�1y9y��Q	9e��~�.|qT.k@�N�f4�"X�|����KɃ�^��8��g0:-��[K�si�L#�"��O�N�{�Yl7�<���?�v�r�(:�/�\�L�EMTQy���� 4�]i�(�L7 d7a���hx�9 ���W��W%̝>EyH;Ҏ��Ҙ~�T&���A��:f�+��˹/��5r'�����W��X��RR!`G�<<��~#�^u`������J��=��腨��9�XA�H�
zE	zBUO:k�<%w)PGn���72�US'����4�15ۑ�݁�_�q�m��|�C3|Mq�hV0�ɷ�)
����t?�$�I��a6\qxyi���T�aI�B��V-��ћ�h�4�4An�`����[;���)��ၥϠNꈌ�"��1m���w�*h+A8�#�bQ<INQ^�c#�qXB��d�64�4+�;*�D�ބ���F��iX�j�<,{�%Ȏ���g\
�[�~hQ0����b�i�6\�+y^nⲼ7Q-Ւa$�Ϟ��`����2��G��^�Z�0�����|��xR\�	�G�ܗ�Ӄ!"[p�A@��Y�rXݝ���P�8|�ǥ�uC'gBH!c+h��o6�l,[� �a�*�Ĕ�� �i*�*n��%ua�rFES�=̀^�j��'�x��_��_DpT ���3о+V��5��Ѣ��&+H�M�ׂ|}2�Z�Ȫ���b�7��N�L`!��Q��Lq�T�z9?B�j�?%cd$ah��Fg��h't҅�#�|4�R�\�LT��V��X[>�c�wЁ�K�K���Xt�臱G��L9��vQ�d��K`[����e9�V�!PR:쾴9DWd��Aq�����?V����n�nD�҆�X�h�Y_��Dn�%aD�C�0!�e'Y��[{o�%u!yo��\U�M#�To���A�b@�؃�����SKӬp"�k>m�6�H4�aPe�1�d�Z-n|�``�;:Fż,W��`��~��A<]�%�"�AH#nA�@?Y�Z\�S]�j` !��Y�7+chrr��Tj����ԓ|?���N����?��X0s�Q\��ɒ�	w,9cԃ�E���Jf�u=�bN�Ĭޔ�w��kx�"3/$��QUQ�1B�0�ڨ'��[m����%�B�ӄ��BS�x+�Ӊ̎��6��@wJ{Ncm�Hg�P뷇���!��OT@ɿ��,�X��HT�z��Ԃ�0�p� �C���1lu�Y��LC#V<j���%X��� �hT�1�n��qPA&4oBG�_��'<'�nu�j�n-8©F�6�R��:� w�V����P�v2L�B�Qj��Ϸ�4�F��ϙ���4�=;p�����9u����kR:J�!i�� ��y4�ď3� VR&W+��(7\)
⤢a^����
�=�Xa�@�"�m���q��հ:�Emb�ԋ!��R���0�.tq!�(�%�����ꋄ�th�@q^�$��MBK7C�P�/�+��?2a�
2@�.�uT2E�)��OZ�:�G"�h���O�.���,���	K��Q���I�Ȯ�߲A��NG�zo;��G#)E����� 	��j$b����"Ø;鬃�9�[�������s���!%^|"��>Z+�)�oA�����`0h�T�����+����l"S[����'�ev!OR��R��v��]ð�f���ԗ�!g�2�K܂�[�̟H[lK��k$���'霐�[Nz�.2qR'N��ĔBT|^�]Ng؁�0b��]�k��\��Y��(��@1�"�3�9�KA"���Y|>������F{�Ჟ+��ԃ�S,_>vJ�x���P{ �(6���H6��Ȥ{&�Q������;MX���g�|����[{�o�1�_�X��7�|���	r�׎)���G]R�GG���������X��"��@�K%=�MkIЬ"j
����}I�p$��=)}�v�|��7D��,�a����baL�����a���� E)����4�:+�I{����"n���g�Qk	�.�a�U7p�K�C�Ik�R6E�����D�d}��m���]����6h��io�)���AȖ�%�������:́h�[<��j�	[1�8���G�~�u��r@Ø����aCG�_���Upu�!�^7���&:>F@yT�8$�I���k?%@p�t���J��>���fh9[�E'� ��Uu8���p��I��Y��ɓ1��
�Ket�# �����1����Ҙ�S{��h����ѓ����θ��*B���+���D�{\�s��Һ�b^��E�Y* V�<cέR�<��dd,q9�I�ǘ���縮Q��������m����_��;������>x���_NsD�ḧhɧ��>��J�O<x�Fh��l����8���{�Et]W>�l�d�Q'��*�5ɤ��q'�0�w�ޱj��W�8�T��'a�R��;/���^�2�(��<�k�C���IP��C��q��a���85�����"[��������K;��Uv��=���Ϸ���_A��Y�耴�-��{03���8tȈl\�ڗ�;�zϞ�[2FWJ�e+u��訩�X��X��c��9cq�#Ѐt0(4�dI����:��a�u�i�C���2i=S>hH������믽�s�����G��T�u��*6�ߺh�/��gg4�j'�B�#� ʝ2�ʁ3���am�/���)SK��A�*�x�����������Vm��9�8�	��oWvq6֦5�/\�(RJ%�|����3h`tB��?�cٲe/�'��;w.B����ß������y��WJ?���Ej0�I_S��MCˆ����i��O<�L�/oQ�J��}���A%�Z��6������-����X���������yc����غm�i�T���%%W����c,_�ڱ�I�I#��+���?[�ֆQ^^�aƲ{R�K��۟�����ͩ�xm|e��\��ҷiVF�����]�x�0���RD�����0p������4���P<�h���'g��TTT������+��vdn�F�?��ڴƊ+��u���{6�yqq���Z�p�����k�0 �[RR�'��v��몪��2�O��hV��k+u]���a,)...�ƽ�o��*]-//�4�KZ�[%%%gfcs֭[W�u����cS4�Z�bŊe����p=�����ٸ���x�4�K[ƛ%%%����ُ���FO���n���0�b�0��������QB�eY"�YUU�@+��m�x�0�?�������o�ˆa��*�|cp�
\�	>?�F�=��ƮX��)]���c�_�|��0�m�16�������SQQ1����V�h4�+k�+W��K&���ceqq1-��s��kM�����8뮽�ھ�ؘ�k׎������0ލF�YɈܬ�]���0/..��{�O>י�yN+�������llNEE�����٭�h4zz6�v�Y]�/����=1p�@N_���˖-��,�W�b��|^66���bRee�V��v4=#k���뗴�Os0z(>��a����(�5��nݺ��n�z�g�e�UZZ���k�u]��3�@ �Ԁ?����(//�4��Z%�KJJ~��7f�ڵӪ���t�]����...�2���c�d���"]]�n��[�n��%kt]�x��?<=`��+~4�1�Y�Z峢�bzee�M�0�\��:g`nI����bN_��p�1�5M��CT���������0V��P�yXƲe˞�,����&�V����5�\��^Ɇn۴i��P(�m�T*�NYYY6�յ�a��y^E!��篺��~4�Ix¶��4z�r������|޲e˖�Y��DjL����Ҭ����� �G��~���k��u(>���X�d�R ��(�|��ʊalذa��͛gAZ:�&5�#G��e�ʲe�^�m�"�G\�OF���� V�\9'�J]o���ܹm�ϖ��e�Y�f͠>�����;��pgհa�f�0V�XQ��'I4k�����,���+'fk�o�sXy����Ζe��i�i���e��nݺm����ܹ�g�i�h��b�f�QG՘��w��A����$Ɇa4���U�=b�Z��6���Q%�H~��8�<�!ڃ�����92f,    IEND�B`�PK   �e�X~��a� ٮ /   images/dc707dc6-8489-41bb-a5bc-77a0670f90d6.png\\\S�� Áh���P%�lٲ�LX��,��
BX�Q���%�A@�� �0Leʎ�gb!��b�����p�=��y�sB��#=�=�{ /��E���-��|��@�W�]~�a�<����7x��粅"������	��Q�K��&�����N
%�����p��I���%e^S����iP��`ȓ��P�ej�l�{�y�o�!O!rݢY��بߚ愳����}���r�Wk괡XY?�q�?�üh���!͵�/V��xt�e~fc��	�O��D�:���s��;%!�E.�o���˘��P\hV��rɘ �;����TS��{k����EA�n�Z��2���|��k$8V�p�N���$&��������Q�9�HO�	��T�{���M�*��o��f���̑��M�<�!�f(nQ����P/ h�fvh̜�,`�*�Kp��e�Wc=W*&���s#�pSx���]jr������Y�]`7�핮��jʿ#˰?!!�\Y0jn��D� ���Ȳ���h��87Mr�q|h㡴@~�K���g
�	��Xy6\���J��ځ�ӏ�u#H�u!�}��K�����%%%v�ou�V'���'���$�
����vv:o��Dz����p��r��gD�*������Tc����u&�17Jw-16������p%�8Ec��Nl�B�{Eُ��^�LG4� �s3�Y&Gބ0�F�٨����?l�HIƾ�䦚 Y��q
؜$ȁ�,S���fDz|�e,�q��傆��Vn����@>$2�r$t-�Q����a��o!KʐĦ���H9�mb�����m�Ž�u_���is��=ۚ����1�r�|ϐ�B-a9~X
j�MD��+	��#ҍ�֘	��1//�����")�	p[�e�5���(ۯ�N3�� d�)T�����ɂ:�x�f�h/G���%�����	L�e���fx{���}~~~��J�1Ε6/c�&�
?LDD�˓��3�{����g?�eB���Qsn>��>�2�+Ȯ�\\�1%^�+���q��>�n���R6��]�]z�}B�u\����uv�Y��H/$�W3�
&d��Z��v���#����ї����k̉�����ڱGw4ʂ��W/��� Ɖ��OP��m�*�E"7f�TU�����a�@���+���=�o�a5sTL̖=),�Ek�k�:V�[o�_�#� �zbўׯ�o��Z�Wud��x��CU/��Z��,L�s�ŉ�kY�����"NN�9�s?���ma�����i�-g�1����H$_g���d#0[��n�����S�Y� ���>snBj���ݗqt2�0�׏�΁J�����7Z�|�2��_���R�t��� p��Sй9;��q`;6����@��VhS���[�0��o��V�e�_|B���l\�Qq���So��D�����[�m�~��B��D,|x*.F�Ƭ_�8��J$�Asp�y�f
<�]U6��Ka����n�����#	,�~��=w'H�g`��w�z�<s��@���Y�Y��F���#����e^w ^*����&���'�
o��$5�8����j�����	^�,-�%z�h���K`�kʋ��Z��**����J`�W	����5��#��i���h!����6Q�#l\Q�¾��%I�>}����t�=y�y��~pyĒ;�H�Xc�u���޽{ͨv! C'����|SE��u@��;�u6.^��~pG��
� �ژ�m�@[�:�������EEE����G������b?�*���������6��7)%�iv֣j�kP~�Ӑ.�Ă���:�tD�B|{B�B��Ǭ�A���*�m^Y	R���_
�~�VP@���1���(g���l����ˤ�E��m6����@��:9߹���п�YL	�i:��fdZ�c�Z-Eջuee�KY]���mUCEUUF�VT����206.���J޲DvM�d�|�v�3l/��i���9����ϴ��Yy���3�;ǲ���9����vnHa��zC���d�?�{w~��|2����r��,D@���ͫ�P�[�kᅠ�,1z3��@Sd��o�<��Z�x��Ey��(韤�����H@n��̮��0���k���TM����PSc���q�h��m(�Y�
-!��a�؄c�o{�����;Ϫ lv�R�
�eXR9N��6��c�ݽ�j�y묬,�/����bF�a���؉����7��Bl=h����>�n��P�J$�\@���P�y�m����_g.$%'7JTc�e�NLִ����������=�g�'?6�L��U��N��=��g�j4B�- %�O��@%���7U+D���oM�"\�"$�p�� {��+#1���G��P������G�8�f^U� �!߆P��ɲ=�Lb�ض�>6ʎ5��-�m��X�7�E��EvQ�K����(�����- E��ռ�*���к�01>�s��� ')���.Nb��̔�98�p@��b���w�X ~*lD���w��-����B�@�=v,Wc��=�M//Y�o�+����R�U���^_�&�}0sD6�h�I#ql]E"k�뾤�bS�4�]��IU�l[�I��^�7���z�5M�뱂��@��l�wTh���8�4i=8�j|�ߛ�8I��
��$�
�}�{<ڄ�o7�C�+S�$�qU#�3�FFF�����r��ၞ�Wz1��c�N�M�cQ����}�".��O����*m��A_��o
GϚ х�ie	+��dH����Q�kE=$��m�2�0E��趖�`;���8�31J���̧(3�ۅ���w���J/�:��K�\��"��PGe�m��=,����Cj!��W�cVXU��L||*�'d@��������Z�2_9�^uj�B�.+��!1���RݡY����)�&)>�B�פ��HkU��k`"�c�/�oS"���ʦ��6C,��x`����vb^�p�`�Q�Ǔ\lsDY�x�,P/}��r�-i���Y���5dx�w8���t���6�#�q�n:��������f�de��=�����Ĥ6)3=A��\&�x(�EE�f�z�����FWG�l�2�����0�㥒���E�i�^��QV^*S� B��Uqк����P�zK�'T��I|���	Tb�&��S����<��51��W�H$5��(�>nV��*
x�Nh��@�/DDD�$n�'5!����<y`3����l/`���O-P�>��-4�һ�e�U|�\�
�-<idd���v�Çw�����<��[��Fj�f��������L��Ӭ�\�:a���E��)hȵ��Չa���J-���`�[0,�)����
\[��&�,5U�����JT��;6�6	)���/�^�� ��gz�s������]��`w
Q���J�����>abA��V���rkʳg�)��:�����wL�^����6�� TT��B�b���9p٫u��ۭl���2��C�uX���_#	���ڴ������c0�N�����{�����J�H�(�aԏ�Ƥ[����ϧ� T���n.I������;�F)rh���bi�
�Cܝ�޽ks��qF�G��W��9�o/�W�Rm�F������'�m�(&�M�h��z�4�0��z�n�<A���(o���]��4����a�<�$@�V ��om���Ź����+X��H��ޜ��P���~P#ʸe 7�v/��k�4Tj��gߝ���8D>a.�`aiY58ƌoP��UO3���f�ח��/K�j�n*�{�� �@Bv��πn����w-9�E�mL����S��0��/.���WN��_��H�&X����Hnz:�:;CσT�����ׯ_����ۧ��V����K�G�۹��K��>-���f懧o�v5�h>@��'3�a������f�ֽk�mv�G<�S>s�С�xĪ���J�Z��M��k𙅅�)����6 s���1K�^��@�z��ʵ�*�P������"7�rͽ����S���q͹!5`*�/Nu�n8�+��4`�0>֤?<������[+�/�?^\{�9�F㾲�N�R�������d��Ҳq}-kS���sֶ&t�ߟ���N rMJM��Q(:]|��}J[��r+�G�	]�E��]\�JlJ����5��2���o+���T���|�j�R��F�Q����v�\x���%cn&�'l�nP܉��X��М`��C�����Mq�ي�@hz�`�KЪ�,��Y�{�III�2̭mlFD����g�*,�3�=3�X�ؠ��i�y��0I�����P�0�v��qUI��.zn�p�f ��a㬉h59�f�~�P�`(�	��D������,J�`Y��G���T �a���c�7NY�{��S�;�e����3lgL� �s{N�>����$�5NN�Y�%@X��E��A�L�`��``` }����?}��xWt,		��8�
`;��	,���NM��W�^��	�`��v_[��xK���Z�
Y����W���eƒ�@�;���+X�\��XfyTX���C�꼩�o�gwk��oS��I�/����ơo��Y��Ü"1�<�"Q���_�|^�����TSZf{K���kEӌ�'�2j-o����������n�9��ھ��(M=�%#T�c��
V��%�!0ܲ�ܜn�*�ӛ�|�`Y��� ֓�Y�?��-S	�t�&r�K11R�Q֊ ���V )P�L`�����tn�O�֏�#K��bmY���Wy��`�:��#֌mpE銰ʗ��1�!'+�i���>��Y��tT���@�`"k[��%�2����0�nG��L \X�x5���u��4�3 V��`h[�V�L�ri�{K�Q~�E�1\�7�LykMU��+ �Z0��tʷg\Ē�ءj}	DrL�45SY��]�i������B�,B5x�s|�����5�!	����jz���?���m������	�X���2�JF�Vh��>���`靵�_X]��f%��}vu��o $�}���6��r5q /,�Fy��N���<a�
���xS�K��4  \�C5��r��/7|f�}�U���ɞz���Z���Y[�]_�ե ��߿GIlMȌ�p@〩L_�0��r��џ<M��}ZV��5RO8�t��.�@�w&E�_X�Z�T�,,\[����@�W���M@稠`Uy���7����h�b�S?��G��B9����~�e7��@�)���������]s��a��Z�u�z�$�{��$3$�����COh����ۦ���i#p���&J�!�;�\���f?i������E��M�gj��7�OH��d�rйN �`?�Z��x�%)[;�n`����O7=����޵��Ngg��_6���~�rq��'&ZӚ@S�N~|�8&�v�'��c]��K�W��1��4r�	�\<7��Z���߯�>��X���IFݯ�mۿ�l�.k;���!	� }	��3�zr�{��]�"p���2X]3����5�N���K��-��ɩ�[k`�Nͬ2�PXo*���r�y��P��M�A�Sk@��=d���*�D.��'{�Hl,��A�� *��.=�zs0̑�e�oQaO2@���U��o�,� N�wG��Q�'V_{s̰�Ƀ���6�⥒ң��������6�@ث����#|pI�e�(��	8k_�g���C-tտ6<�'�W_�p�ڡ���YAM��&�jSب��}�_J烜��X���l���S�n�%� bSk�P�1ߟ �he��X����<��7? ա�8��J���X����k��<^㲭i"��۱���S�A�M�T#rrr�D ?ы�\g~�(QQ�fV��O%���,6腟g��K`��<���s90���4X?�B=����/,���~�2y�a�[�� /Wל���!UY6y~ڴ���4$�J������u�g���W�}�8Q;^rݹ���%ǟoO�z���U�}�:[$�p���y쓣<��bmi ��������?�m�-O+�T�X�������u�2�xs`p?@�C �c��B�R�m`��0<ˏs,O�V�x�$�C����c�'V��[S-��K3�k?>�Q#ǧh��8~qnC6�������\K2�L�h��X��ꇶ�˓�C��Z�ִ-��@�Z�E�Y�v�5��1�ָ+��-��ָ����%��E�s��&��s/��� �mqwb�X�����|a�~ds�g{�B�DA{Q�Sqc������D�]���Z��,�)��y�X�O�-��<�շ$׏�i5��ʡ`,\�87�Z���n��`j�\�N��.��o���E�����{�ID�$6��!�?/"6{���a0Y�*�v��_:��ء���~�.��۠f��a�c���B5�:��ڶd� m��V�d������/��R�й	�����/P[uC걣���\Ǣ�H6�e�ϫ�J�PuףF�(#Fk�l��� ca��/x�����&�=��r���3�!uQ���{����J�>Q�ġz�h���I_+�1�L���C
�A�h��C��\m�&�O�j��P'�uE��)��a���������˾�ޡ��r��SbƢQ2�1S��ݐs�;n��D�m�Nw2G�Y�!ayO�O����dY,C~U��!z[��K�����p�<ۋ�|ܯ+��0�gϨ��m�az�	���5�{�RMY� �$�lz`tr0�f�� �G�v�V����:�_���Ƚ]�wC
������r��T^n�Q'���n-�xM�$�����q>!^�h9Q��c�@nא
�Ճl�n�_D�/�����g�k�a�2b��b\�4� �?�e�N맃E�D+����0�j3F��
vz�A*_���p�\�y�;o2nt��.x�9�qAa���}�1��J��
u����$��&ɾ?q�h���}Mؔ���2�����۬$j�_�[��A(�;,��+��I�7��A�Y��m���++�O��,�$�d�����ȡUFH��(�S��:U���w������!0��FͻL�5�=�g��vx^_�Jv���>e�b��Lg�V<=_�8��h��>y�0���61���j�O_��������@�X�p�:I�2�qm�/�}��RT`z7���[�a��V�bSL6��ˆҷ8��7�WUH�]t�PI��)c�1ùw}`��[��9j�:@����1h����[3d�����{"4c2/n�j��;�aw�L,a�p�`����y��C��c�kT$y��3�����8�:jR��e�	��g����`t9
׵=T��
H�w⨟(3֧��������Ĵ�1�Q&�m������߁sHw�7��1�	mK�m^����Z��rA�y��+H�b��j,NO�n�"Į�HJ����s�d��!}/��6�Š_@u��4 ��w��(μ�4��Ѻ�#*���t,0vRd�8ǗC7!�v��>�S7�ǤʑA\I�3?Y���H��U�y�&�v� ʴ�i[bp����;�E:��:Z#&��a�ua�W1ߒ��HUY����ˁb��D8�_��W��e�����eGL8_%���ȉ1�$oWu;B
�?�a��tT���Xm���ޮ��:K�pg�����$̺�w���!��vz<�:KΎE+��j����qj�}J;J8Y�r����B��t��:BS߼��?_�Jt�vMtGF,�*,C�p�G$]�	)���ȵH�͟�O����!KOz�ۤ�Wwzn_)W?(�OG��>-I{�N�)U:�a���;i�l�jw^�/�VCA�]��%�W�g ��/ӟB3��7`DsL�$9�U���er���4`փ1&��Q旗�<$�1�3��`.\e(��:��*���C���3��ѧ���"����N���=؍��%κ��
+R��8��čA�.���2�p8�Zo��tO�v�h. =X��	;�^X������`��G��v�����e�3&F@1���`�������A��;D��0m$�0������/�z�}��&���60յ�� o�v�O�*%�A��ݳ�bz��K�v^a#e2h�8j�O��`+��9�v����O�&� ���T� oA��&G 7;����ϒ�H���ə�Ab_@̏�h����J���/�R 4lg>����Xкщ���̋0KV���.�b�����OF/z��B�]��#v^��1�3�8N�N���i^������xЭ2��dE�+�v����@ƨ�(����H����L>����g9W�1�=��i�Ϯ��o�-M2��L�+uw�6bGj�� ���g!�۽���N�����#��h���!Q�!��w:'�ea��Gb�YP<���W���<���j'���@��c\��uŚ_ND(_�y�[&�O�b֯��p�9���-���´�1�7`�]'x"Rv"P�N(,�d�%��,9 ����(G �XM3�\�����H�;X���Z�ť����>l�W���y���?+͇^��)χ��?y�9}e�yZ�X��$��c�i� �S��Mi�}6~�A�)�����qh����!I)���	�1���9,L�<lL�@"��8�~Q� )vdd�*��2k�Aɀ�p��H��SG�����!���p�M�1��Q,SHCl�P��x��^�tG��_�6��5Ka�b��`� d���/���y�L
,P���0X��N�K�bg�u�B��Ǝ��D�������G�Mc+݅����8#�o�&�25D������jV~b�u�3?y��������$kY��y(��G�01����u���hA�0~l�����ql�ߤMݑ9��2$"�s�h�]N?���D���Z�#��������D��k�:�8j�yۏm��([y�d������]��z�����ioxԐ��D�6/aj�Dk�� �_f�/SFM���l��s	�ߐ�C	�C��v����V���2��5��S�|�����XX5tNGŮ��SE �O[mC5=����	1�n�G&�ô�{���WN� ����'$���o)?�QXH82y���g_k��+��vG�������߂{�=-/���fk<>�d�Obnn!_}����o��r���-�rl�����d��p[O
���kz�����P�W�/\�-�=~��4r�=��_������?�|y�TJb.��H�p�)k�z���i� �=Pأ�l�f�����(ͷ��)p�?j���{��۰<�j����ϡ��צ�g0������\��
� �|��a�b0��\�;,ƕ��8�s��'7��szr�ߞ�M6��>*�6� B��<��9i�N�}��u�	�%�ﮦ���%Cs���$�Qҧ��jm(&Ց�L٩fl=l���8��;ҾlMi����W�M���E+�zp���� �?2��摕2�����[-�Ӯ�_����B�{���W]}����E�H��e{���k��>5]�i�W*>��H�P��ݭ�G)TD>c��R*�����#�ɐ�~A�Wr�͸�x�_t���T4�/�׈v�����Ԁ)7�Lo唏8-"?Xͩ����o���k�w�'�y$2�����,�����Z�b�ٌ%ņ:��s�N�g�)Ƒ����(1�M��ɘ���Z�q�q�EA��{�a�}Y��S>�+}ͷTB�(��T��"�&�Ά��}6��>�}�;�JH}�[{�(�ϣ���%���[��!v�j��(��Y��__t?��;Xȱ"wp�+���3����kֶ0Bm�0����1���q2���@�����I��g3�"�^�NTŝ��������0ب���U�0D���7���aK�F�罹����g�+5j^��q=|;G�= -{�BY"͜B�ή%�,����^��o�l��I��HF2��-1˭�]����=�o����}D}7�����a�߹D0�WЍ�0ą��%F�9�2�$�ך�:h|%�y2������rYHJ����ڌ�)�鄲�|)c�쳻6�8'p!q[V׃=E�;L��K�Hi����Y�G���:��[^G#Z!)���Z�@8lE �^��r��ݼ�C��4}U@#H��*���Щ���W �"H���v+`�T"���/�3���8H D���p���ri�-h����A�� ��4<�X���k�0���u��A�]�<>J�����3ag'2��� �����V>����߯��m�&)�Q�H��r�L��� �g��;=�РS,S^��8Sg�u�G&B
 ��o�d[^�=�+�[z =��{���e�ο�Wj��fa%�>���ɴ��ڜ��i�*zC���Þ�x���Y�o�75&����];�:�
�ŵ.MS<�ͻ��5Lh��M�vi>N��ﲽ J��O�+[�¢θ�*�7�z���yv�%��a����Ӝ�P��Ϻؔ5����~��MDɽ!� ��0����~li���u	Z�AmȀ�sV_���q^���O����N��J3���#��m�؊2�!���FA�n>��N���df�)|z�<�>>��$��"rO���M%���&s���32�1�=Ј�����Os׿���v�ushD4�x<����H����:������-m�S-/M�/I�
�szq���f�@�M��X���bczg^C�:��/�����ʮ�]�f��0����U�	vmCѼU���D�U�� �v�2~��O�ē��ǡ��.���(銎�����hкL�_�U�်�G����^Q�O��(�pT�����]rf�	��Y�)CG���\�MON�&��U�Q=��ݯ_�C���>�.�p5)=�98X}N�󮺺z��R�vF�nC���U�lՀk��I��p�u7�u� ���FS_V�!Ô��so>==ݰ�Z��9��E����b�F��<�%���Q�W�W���f֝NlRް�E��.��ux����o�ᝨ�E-���o8-� ���t"~?���jDJ�D�qU����'������+���#0�3ٜ��zz޼'ѯ�|_�H��uN�������T���kB�(�PiӕCU��3)_ߺ��^��93���X����ٳ˞�����4�k�}����!ct�����1]�/6�a)��R��~�ʸw`��x���'/���.�����xe�n�miӓ�'999Y�$����7�/!6������N��8� !��̤�%�u�����y^�6��YNWE� v������jЎS8���dwGxCPl�Ӿ�˖����̳�u��8�3�[y��Ŵ�͛|��G�$��W�X��,�����ҥc�G�ʌѱ$F��F��,���ʙx�!36�D��gm>�t>���~��bFb)Ԇ}�kY����H +K�ԇ?���@%�@������D����-h��E�>��psE���"1ؒ��v+�����	�,�_`��/М!��h[5W�=x~��	�Oќ$��l�9�:"�Exl\���^���kV���o��l��:���y��8�G搯���3�9� U>W�٘�'#�>/>I��2��{>T��I��!�aBV�c�}��|�PݯIG�Q�Hk��Ʃx���=����h��������Q޷N�m�i�}���~��Ec5��ƍ��"R�?�˶����uO5�@li�4��oyL�Dʦ�vJK����9nF�[��{e)ڕ��������Y��3q]ۺN���͹�WD��
����X��̺W����լ�
�{�����+����3�cqM�b�q�[�o�}B��Ç�}N�&b�����7�Ż��8�+J@+��g�� l�s<�}y�=�Ϸf*�;:�<1�~?�*�)��$��,��(l��P=6�<n�kk��<	.
G}+�=�Μa}L�]���ށd1�!��n�>̪�s���>o��2h$MD���Dj�׾)	�k��o��?)�$Bd-�?ݢWg@b.�t�|�!:�t�	t*��L��s���Q��$f�79��&B��$&�4�6*�uZp*^`�M��)��aa�	�Esqǟ���β�J�vp�T!o��#�'h!����ğ�$��]���М��"?��-��k9`���q�����BeG�K+_(��8�����cxY>��1�O���Op ٘�W�b�PS���Vz����U�oj��uU�.�c4���sw{.ތN	��m$]����r�~�z�L����|�uM�e��u*��<O������L��11�H�3A�mUcz���HʎH����co��m�8�3��.�>{i��/�p���7��Կ�DL]�EtP]]$i���Pl`ĂA�u�����ԗOE\OJ\r�nN�byZB����\����Z��CS��sKh��9l���3�^jn�?�\���,#�Dz�#��Z`�'nPBI�S�K�'dRo�l��j`I-X�j�7�3>�[_ooR�n"ayI~.�%�����RNhe�3$@`�O�k�Z4/r gyt%Dr�Wf���׻(�,�VMryqE�&�}�{(����	����' B��^\��{8YH�[�$_Hf�{?��c�R�kL������0�F'��s������NIF���\{�����<�˖}�s��U��)W�<-��#��&@�$G(��܍��DP�B[��<��@J]{��T�B����ڢ�#83�镴U�tٷ��"ü�h�ZyCv=fӈ�5M���hő�ˋ���mӋ���/:uޓ+"2��PP6[ͅc[8�e�����>�~�������δ>>ӢEP2��|�7�w�k�
�}ө�y�p,���S�<����R��ܛj������w��_�T�B6�tH鷿[�XEx_\yų%UN��]� guv�_���4C��φ��o��Lm��U�)�@�D��d+x%������b��"@�lv�����IR�;d��!���^�����In�B��4i��S�6w3���x#����U�OTG0�Wწ��;88H�U.(U��k��搸�Ǟ�����l���k��sY؄@�1�*�J�R��^�"�/���2��:����5��p؇�M;(kH�������d^���/b0ݙs?Z<�Ry- ���������Ч�����Qw��Q���ޙV����I5$������+�%g�S�b���n��~�qe�(淞�*�ȗ,��!;R�ҿێȕHl206�XX 8Q���1��c�T5nӡ���ȦR�*��SӔj����:0����hI��2$K��$�N���>t��)��Sq����۷��={��u�q�)��~��%������=1��)�I��xS� G�-�?��pN��Ԗ�����4���,
��-�r�1=u�g���lC�}��E�u�ԃ�G7��i27��cҎ�{��Y���Q��&̚kW��ێ)�4]��E�{`Z=ǖ�{�7�NI��X2�·��D��t<H����%v�~�^�����S������ �X�v!4�T����c�#���4�-c�j��3�ʗ�bO֯<.��dT�DW�h�ة2��Ə
g�����=|��|�����l��|Y111A���n{�B�ȱc����Wz1b��j&��"H������,մ��`���Q���6B
�t���Kk;K#'9x}�Ћ�/�M�t��/��I�N	��xC&�Aȼ䪲��zZ��Vr��7����u�h��n����(������G���z=ο8geulnn��W]�>���422b`d���+27�,��I�5�-��8��[��K�8z�͹�-Ȱ��+�w�mS��l>ϣ*G]���-LNM��l�����L��Ż�����}�J�Q�n���:�d8j(�C�c��P����-��-=�% ���<YAJ�t7�݇V|��V{���߄)=�5 ���[8���|����]��G��Y���@���'�kJ��텅���r�t�(��[�| �
��:}j=��e��$�;��g&ք�[��?*
Cph�UK�UK�j.㯜��b֎r�7���}!Dp��
�R6O7�M�k �b�Z��9���1�{1��	���@*gخ
Π���3�}�iڔ����h/ |`S�,�o��L(][v��;8�J.�e�ށ��1_;�1��f�F��6Θ#����&�氯^�����t\#�qQ�|�8���Z�.������R.?�vY,V�7M�d|��S�5�C�M2^cb0���Gu_����d�Ӈ��F"�bccn�K|���_��f�U�V%E4�M�� �"��$������6VI1���|w�Zk��`Ւ ��Ix�F�#�}���m竾wa\����ڃ޵�y�!���dn �-�ڴ����@��=�p��al�n�������O��R(NO����[���=
m,SM�>���ܯ���.Z׍��:<q)o$�8�PTW_m?2��j'�y:;;�}�c���7_(o�z}2gI��s��Z�ZK�|�"�|(�^:�to�+�LK�?��tlJ�)0*<�l�eڻ�y�Xd�35Y�J~Rc� ��~Z�U��(o4lA5���\��G��)��$cX
!�����W���z���͑�G�U�%e����[+�ؔ%�.�}��X������VO�-�N6Q$�=�0�Qݩ��乸��;������� ���@TҨPu]к%vU�e s�I�p?�7Y&�*%��fL8 �e�^�6�����o�2��=I�Mxw<�7&��{��8Bҕ���^4�����<���/F3�8[;i��t�8k��P���P�K�����-����ص�<׿V�;{��; ��y^�՛�Gss	�U��MdM0�{����u�|��<�;v>�=�Wy��,����oyY[�n1uݼ�v�Y��	`��uCa�:R e�t��X�M���\Ȗw1�&6���[�����|fT)�JV��z�6΅��̱���%_��\���s�Yw�$����sz�������;R�UKi{� ���4Dt'����� ;(���*# ������FMf��o�z�0=���wz���}x��`���w[�|��xOrƥ������0��5s��D�1���rϦ����8��zR�⍺=���~f���[��� 5Wx���Ytmk)A���wK>���V3W�O|f$L�XD[9�������{��l^uҋT�Ƚ�CH���k�B؈Ɂ��.A��L�>bhH�Xl��]��ݟyް��D��O�(�^�Y��~�]���c���֯��%��e ����{翼Ɉ�/FQm5����'�$�``���1�ɽ��|�,�t�@������9�\g���h[� ��d���3k�yJ��D�"N���u��$+ל�T���LF��I3	�Ћ2\\�{i-ۣ��9��7�	��-ة�����t�q�ri
]�"A�ȹ&�c���`���`胭#=��O���T�=���0����M��#:)dǰ[���#�V�T>a~�Ź�#��m�)�	�{-O�ݬl�!�0��R,�N���ʙ+��`��w;t��.[���ϯ�h*(���((�}rr2tI�*�@̯�����JG};�����>�M#\�s�p��m��7 �-}?��vgؽFtm���D�쒋�3��ߢ*�Gt�����g�}��_��lՃ�=��Z�.��}�ֆ+����ߏ��mgv����7F�\H�@���n�{-05�N���I<��D�q8�7چj��r���1�9tD�s@��@�����q��SXӧ�i�H?+�~�����T��������<�J�"sM�;Q�|��YY�#d��.`������9�����`m�*g��ܑ9�UZw}�>���][0ӽ�yW�J��ִZ�u�<jӘ�o�.I�n�y*#l�<�&�V����9�L������1���.������7j N[�S��@��myfw��J�G�@���EF#�3����w�ҋ\{��5�J)|��;��'����K5�W��4��: j������F��	�I�?�jP��I�3yb��i����=`����/�>� ����=N��`��=ϓ-�4�����g먬��43�8ywA�뵳o��C��g@��� ��5ꔼK����8��qV�����o߾������>D5t�����R�e�Z����3���kI�sW��Ԛ�m\S`�Oف�(���1qq�CFY;t?ۖh�-����	B6q�ޑ��˨�vZ����S�G�� 3�TVF,�r:�1Q�������]����O��X�,�,�o��aٮ�ȇ����V�5]^�1q���!2=��S�<�z��m��jz����>��~� �G�qh>�u���}�j8�q	��2Qb��x�����^�c	�f\�&���lPI~!)O��m�~lW�KL��� d����g���\�����Mw��Qr,z�j���5�X�QAAvʿi.u�H���+)��� (J��CL��h�摊��59���S�@��000������]�wo��^�=���<�0�4hF�U�IѶ��n�6-�?��8��W�_7���D"l>��z_���XZZ�q�gb�y������=�v�c�Ho�J)%��9��$�?~�/�XDƮ�X9}�	�]@����.�����xY����r-[�eB�d�ۍ_��+F��]N:q"���o������ֲz�a��?�����Mֲ���U%�M���t�*!H<���ag�  A���ޒSS�ǚ�Xᣇ�lu!�.��N�*$5OQ�J�V8>�es����v�j��< �E8/9LA��-��>V!��M�~��߻v�ĵ�$��rv�r��$ Odyy9hy#̗�/NF�������Ϯ|��t�3 J<"�f竾�	�a��+1 {��oY?�$��$�Ν/u|�����U����}��0�����׾���u);U�%�)*::L�~�ڞ�Jw�zj?��Xc��p����S��9oo9�ȰT�|��Zeo�����%�d�qL�B�w�b��sm=�:�a��JX�;ݞXz�3{#�Zs::: *|F?�>����8��7h�ug��Yڥ�#�p�ͫz��hh�=����-rh�:����wU.~qcmMp��8�E�D]�А���m�?Y��Xp��M@C�p/�cmPd��-;-�bd�Y��rH���+��[��R8d�g��YB��$[8[�&�~�2�xN��x��N�<�ԇ�C��{}y�, t��ݞ��"�HK���嘪�h�{��?R��>>O��U���LLL@n  ZsL����I�N���J`�VI��u|����ś�}��|��~��3y����4}w<������HV��Q�){o�P�̮d�ۑU$:V�)#d��1�DI����>N�ؿ�����q�sw�u����9����K��۷o+�c����jxԝ���^��j���mO7�*��&Db}	A� ��'���l����Ȯ��Ȇ�_�i��9��	��.�7��H��h���R��ǌY��b@��zM4��Rʬ�S�&:�:���)��qb��O��Ƀ��>�d�r���3_4~��
���J�j
�
�7b=$��ĥ^�: ��,R-�S�9�+]6�s�0}o�h���r���g��X�+�5D@"&���)���ʎ$�����4��G��z�w��"d_�~M�r�xH"Le*���Y��[���-�Ժ�x��Kz��ri���������{.�Ba�7R�⩣u<u6���7���ɸ��No��6��0�0�<�X��MZ>�a�(
��Ȋ��2������N����P̼;�c��a�o��/��HXy)y|s���=�d��	�VU�K��X��-xWX3i C	m��i$	PW��dI�CF�F@����Y	�}�F%���:Н�*���&�m����|-�~�a�g�B �=�2}}`���M�^����0Raa�=Ț�pl��WͭF�8�ח��lh���h�Z��R�؉dg��S��]}}u�)r���e�s������6�!�M�f��ք�T��X���0.@z�`����1���0v�ҵ�2���T����j˶����SW���"N��P���S��A�k��z������;��謽��e�)��
v��$��-^",nG��TK�Dw��8ϝ��M?L<���A@*i��=1f%��%r�]W��@Zk�G
�:���F>�=K�!�J,t�.SN���:��U-��#��/:�F�n_�񵛮'N�ɱ���V1�P�Y�iW�۩��_Қ86A�\.'�=xU! ��N����g\��I���T��:�:�ם��_�#� P�e%�`���A�?Ra�3�P�- h�4d��Fg�KS�y��^j�#19��=�R���8�d� ���{^�m_��3�$�c�|�zu��7���C�*wBBT�aůݰ�21XY=NV�\�L��%Aqpi�gV���'�n�"vK�����嵵��ű�z޿��4�W~�jjf�d�l��m��7�E|��0� m<<*l�h#�,�kkS������E��ݱ�P�nn������7�sQ�(��Z�ݥ�\�TV����Ѕ���((*���<j�a߲l�p3|
4�ň������=&��yyy_fY�9>����<<��9kSO�|i�%�����w�G�K_;��f�L)b���Z-������c"bq��e�Qܐ]�-�!����ֹ�L�α:�%k
�O�kg��K��XX@�O�\�=8hȚ7|�R�htՌ�H�)����w=}(�G�>�V�;A�����w����bꕦ�����K[A���s��!?ޤ��)Y-H�l/w)=F��B��k�����;=�cn����N@���
�̋_jkISk%�Y�ѹ���7Qi���:1���Η��T<?{E���U����٢��v����Dh� ��oݙ�+�T<�������BXbB<@#�LG�$
�|�yt��8��j?1�e|Z@��~����CK�Zh���t_jl���т���[5u=0 �����h�usVK˭1s�5g��x���c�����\�2�ՒH�������w������^��~���X�������TknPbecc�l#v�a��$��7���1�� A%����C<^���	X����\dGG��u=��M{��^�&_�yQ��y�e�`ޥ���qmZ_Ta��zp��2��{s���A=��Y����%���Ö�/NB󌽩�i�K�&�P�Y�3ƹ���4�C1�W�!2�ٚ�T�K-;��x�qq��x���Qw�4������hσT/��@�G�8rz#K���qo���o��A��8���{�v�LF�"�'����]Avtv�J���y����.��H���x���(٢�M%�[�F��E���$+5�΅��kK-h&��V|�����+�R_m�i�)Nω���(̉����>>�<0 ��ׁ��P�(_���rTn�9�J2�IDs1��'6A�N���iLqޫׯ����B��z֝���.��7@��݋���x-y<<�D�kg�Z�}UUb��	�k�����	8�V\H��OLgI5hb�L�Qw`�j���P0�6��c$��7[���Ν?��l�����-%6�8�I�a��	,'[��h���\����/r�ξY����^�SZ_���+�+�D�ٲ�$�K������3��:D���k���?���g{.M���z0&���rO_��$�A+�������)���h�1��0ڲ�G8�n�@����!CP�P( #��R�=��b���y\S9^�~�b�Y��߁&T'�|�G�,z�I�f��Y(��v-��������u��g�4�C���Z��r"��g� �W�V�N���Ъ:��gF�-�~�8��;����z���Jի�ݻv�͠�;���k��H�1��~�{
�p����h���[�-��tQ�w���R��?���vv��|�6Q,�ÿ�����D�7�:w�}��͸흢p�K 
��G�ݎc���4W�t�=���w�Q�P����
���X����ͯ��s8X��B��>�F�����jdC�eb�\]4�ąN��/��Y��`*�s���m�EqR�R��2��f�(4�U\���	P�����x��GQ�
E�m�]D�=��ڀؽ���'i�+��tޙ���ӌ�;��TKK}�����\��gJ��\ZhGy��mv��S�jyd Sd��C�~��!%������.V)��HJ��F�����<.H��z������7��s�^�*�G 9/D���lv<�.�龹�~w���=z���6���%=B����0ۅ��Ҏ��{@��j��慆Z�Ǯ����j�v
Vy׹�>'��5x�EZ�	k�����ޘ�{�T��9���K �G�L�՟RY�
�D4z*4X��xj�5(����7Co��Ih�JN�o��*�����_� ~�R=�e<,�,݃'v`�LB��9����,���-��M���qj ^�~�/������S����?y;J������=&�me�
+������s��k�4�j�f���=������T��t����??���.Pϼ��ԏsZ�b��=��T�՛pZ����*�>��j��܂H�FMo�/��I,j�B�D���"̓BִY���yd�ʛ!ĩ�9���C������cT����⧶8#&�r�P������ڰS�-Y\s�O5q����Ai��$���jn�0�bTl�����ϩ��v��+�nn��3z��/���r-�6ȸ���}�x����꡻�����nMMM�-k���U�<@D��|�r�2w�!lܜS-f;E'����y@���:�R���q��ϯzt�B	L�i&&��8Y��^�]�T'p��^�z��$t��J�=X[�s; ���H�����F'5��B��Ȳ���S�Uq��P�\N�Q٥�TǗ�[������>y�����~��,�������2�wr��/Ma�9_�[���|P�X8-B:lF��_[�ia)'�IVZ��v�nms���� �7��/���2�y@�VTTdV�����s��bU�M��]��c!nݔ �E��5I�^z�R�K�.b��TC"��R+ɺL_]�h�z�+m�w���3���������9 ��9�o�d��+��� �쐏�����D-����G�N�k�V�P��~� K�p��`��l^0ٞ���%i��l�Q���Q�Yyi���mMf��{yAA���w�R�4i��bg�����n��)��q�����-е}'�I�aJ���昹k]��\4B��-�x��ew��?o�w"B쮉	'H�'@m�y�&m�l����~\!�V�������=Y(;w7&��D`Y�T4֎�Dc����!}[Wr���,�>O����ɣs�S���(���ۦȦ>#��:Ew�~�y��g��jڼl"27r\�󗏿*�6.��p?�"��(�,�[�6�d=���P������h4pN��!�y�����-��,�L��`�6�_�֋f��r
��Y�*q��/���(wW4�����&�B�Ȳ0k��шL�ٿfK7�*oߦ���u���B������@�L�_�޽~:�z^l����P��59� ]F,<�C0Rzi��`,&���x"r(���L�A	�	T�5 A��f�#�M�+ܬX�v��x��y)�����X��y�yX6MJ�ib��6L�<���d��ރ�0	Z���b!;���6���ϻ5F^͟�A�GEG��U�n�	r����oR6�ƪ��LD�`>(���b��w���II�m�����鯘Ab@���s]x`�rb�^ʂ�|V~u�� L��z���V����x�Y�����V|\��NP�+sm��]00��J�E�R,AP�(�]�=4@b��&t֒Pj���8^�ؐ"K6n5��_%;��+�LA,������Ä�8A�6iF���R�K����5P�1@��3�o��݌ƙ�B)�ϐ��>Qo@�d�����{CY�+G=�[�GLAAa��حE��Rc��T}
]�VQ6 ���ߚ;�s-���y5;��{�/��E���Q��h�� $�p�f3�jk�����E����k� 9`p��:��$l@4d�is�2���X&>9w����徔1A���ǯ�#�8?�a`^K�2.�i���@ �6�p5�j�bNOM�|�9�7�P��Y��g��8�ݍꍐN/ᘻ�W�_RR��<AE�N8�l�1fn�oj�o)�c#��'���?g<}���dߠ%B�n�[���W��	�Ф�6i�,/�*w����U��/��6CEF�q�3j]\�Ҍ��ܪՕSf��`�нN�� �F�ޫl666�UC2Z��o�˛�<���ߺRµ��� tg��5��<'�I��Qq�#�`P*m����M[�X �� r�V� )�O������l�KuMM����+3=!@B�Q�S.�q�|��'R"(g�Q��i*��;��;l�K8��������g?EtТ|s-:a���K�*��xU��V�0�0���gǬ"`�и����a���ճ�E������)�,S��Iڭնxg*���?4���� �f���Sw��6�~V#Q����VM��,�vq�|t8����<%`a�X��G(�鬓��2�Ɋx��v}ح4�yt�XvO6S%�ӒJJ���[v�X����S1pC�@�K�9����୏VD#
���߾�������C�7Xl:x����9����1��/��28�u�Ctnۂ��P'[`k6�{S�hw!�h����l��YE�C��HލB�˅�3�TH�g^��cC���7���~�8�n��îJ�8�i�ޝ�$�Ey�R��,�@��y����&�����
:쪒�����qR"�^y�M&YN8����4�q͏C��]n![94�d���q5>����V����^�<B��2 ~���*��zWW�J��ZN�����p�� �����KKK�;��Vl׹a���s�YYYP�@&^�o��Ѻ�]����ޫ��=����4QWW!y�Z9��A��uS �#�R 1��o�����9����CIR�{`��f�4�l�6��R'��l�^v�Q�^E8�k���X�1Ԧ��=<,hx�ʽc���A�����P�jk�1��ڃ�A�<������{�1��*,���gs�������ttt�z�ѥ΢�9�������ſQf�[�n�黻>*@����@�����=9>�.�~��W���i7xh�흝L�*�4 �/6�Һ�0���ϗ/2�%fmEF�:��z�\��ϼ��}/n꧳�������T6�����;N 1����??h�6�.�2O-�Qy�ʃC�*F>O�|����º��K-�g�R��	9Gv|(R�2�!F�#�:��2{ՓrS��aS���I(p dr������Z�󎊊����d�kn�����72y�t!�$���1w�B���w�IF�l4�j/zӹ�����)u+h	��z�X����� �`m��/�+���g�.�R%�]�H�������ۺ���ve�i��jӏ���loKὸ���"z�L�"���A������|�H��.��1�}��Y �yݙ,2݁���4̂tvK���� A"4���%y%��v�}|4ʗb&���Qh�o7�����~ỤJ
K��A"7��#D�_ju��h*�>kʤ��[� ���ci����ԤRM/���ա��Lȕ������s 9�a� ��6���f�Loۼ�*?�Dg	�c*�I���I�_3�6�Ղ�������s��m��h6=w���u ���܇V�a���X͝x>���B����@���ܢ�����B�5�2􈑜�:�y�?�43y�/�\��<����!	d��ϫ�Nc?PXĊR���)� �O������T�׳��ӌ���+���\RbƄk�"�"(˟��K��E����eQ��I�
i�?tq�C)B�;���uo����d�O�2���LSts��ؙ*Q�E��W�?��Tf;�W: ��q��Xl}=+={$˃*;Fȝ�*S"��x��.������XkH�픗�w&�J ��x���g���f)��a$�wG��>��A��^�}�|��"#��z>�LW%���$.H���S�cFӤ����]�1�on�p�9*ZJ��6�/7:��}��HO��Q�^o����R�l�[���v)��g��6d�0vO��F�[}y�;�F��C��A�s"�l����K�v�f���{v���h���K���v�C����\�}��F�bI���f%�:�{{�
�L%Ʊ>�{�C�}|R޽{�.�E�ͬ�=�Ī��Ē��e���u-��1��nX�Q��]�h�}�؛Y��|[v!����Q�ˊ���g��:�#jN.Z����ᣒi������^�����9(ం���\��4:'�0���,�~�{��@�m'GV����׹s���?d*���q)>�2
!	�e���ܳ���A��;��Ж[���!K���᥈B=���ez~�z2~.%�y���X�������	=	~g���k'�r(y��VLH����ݠg�����d�O <�Y~J�n��W(��h���v��=�ⶎ�+�p"C`+�G�vy�k

�dn>>�Ý?~�}��5M�[�|��ș���Xrh��$�-��6H�0�4��s||��]Ĝ�_6�|?�D��5G�DV�%��&}�S�D����ZtDY�*�ߤ�x��g�T��SXk�DL�6���9p���v6�������4�$��,�-�]���E,C�(��c�J��u9Taߓ�'H*o[$��P�f�`f�{�@�B�T��NT�j��:oN7Bk0�N�	=����S�ר��[�� �X.�.�:��r�f)K����G���p����ǖ�s���|�k-�ئ���P�_�ʀ	�
?�T�}��%���Gm#��^W4�j�e� u��=��5h��h.5].�条�df��������!@���RC�$�Chjv�
�o�>��P�n��s+��3D������²��Q��!y�2��sՙ�H�TYp��LΌ�g+e���;�+#�i䨕8=I~pBz�1���Y�}��tû���G��$��z���I{zv�:��&zE��h��$���-Ռ���x5��	����
���QQЉ&ҝ�x���W=0���nԝ�ݪ����,��Ʋ<��i�#��B�����[|^ԃ�����<ЈGi:P� ��q���{�$oܨ"��l��9������(^�nrO3�hyKRA��tc��W�w*�R"��@B�EY6�Ю�N��,n��H������A�/���(�r	if�r�P�X����Zw��6�p`�j�*#	a�S�3��N�ц��X/	��?d�CʒC�no�/G-/�"��"���Z�z�$q��+��~=yv+Q�&�=�9 -��s�C����wC��0��c?�Y1��Ձh�����i�c>^Պ\#�Ta3����"3��v|oCd,+�@D�����Tn^����n����Cw�CS���Uk?Gߴ������EN�@Z�ﹲ�(�z��:u:�� �NA�js�q�F�@ΐ����Y�E����8��0����y�UiJ&III}¢���իW�!䝯�}���m�#?�$�oA��	�F��z�̴���z��(����������&���N�s����M�5j^Ck�>��]�M��;���E�~}~��m�Yh?�#�7�%�;qU����g�է!h<d���N7��u��p��,�*mCł���	E�]���'j��{7胸0p�j��8�iEI��w�E�K��Y�7v	f%)��֟a�7o� �g��"�|��Y��7^�<./_h�%����L#p�_�Y�g0�lfG��l׌+�G�{�	"��u����q�-Є6�sr|�ZX�Ub[8*{,�~Be�� 
*֞�+x�N<�xL��Jx�@�����?ڭ�qZp{�D�籋�C���/\�����NY�掣�K��x���zү�X��Ú�u���%)y��[>?j,Y+|NԮ1c�.;��������j���y �9&|~���:wkѯ_�����z�0;�Uyu��4C����٥h&�9`��xAe4�m��/?�Z�C�����tm�]�J��i�mt��{�3� �o��h9׶�Z�9��H֪��l��s��#��"Q��B3w��2Y�xH����0J�K1�����׼�ѫ�F� e��1e�����W�����.RO���G���؞SRQ�k#M ���|�s|�s��p���jzSJ���0��T�����2��ow��H���?�(�1�.p>����KX�J�!�r��D��ۑ�r�?-�l�0K1�o�*t�[��|����&_����Fq�/.��k��g�U��Z�M�������H�r������A�m�=��� �x��$+�]�
�v���XQ$�
�xLSN2Of�b�|)g�����{���ljt�������d�YI�#[%`]�:��S�F��~��p��y=9��#�n��Wh~2��
$ag����hĭv&@^�"��g����b�&bd�͖q;2����0Y���%=H�v����|�G
�a��|W+���r�>�)3.s���{��_���>f����Ĺ�K����˨L5n�*X!�Sr���y���\�7����!���ͨ5�5��}��z|<ʍ��Â��E/٠��V�%����8��"�$$��{���x;8|�8�ݕ���-Z��c?�����V���K����e��\�����bh�X�b':n��{���@�C���=O�|�G[b�0�LM[�͉�u�"��缊>\��9�q��s�1��ZI������֤4\"
G��g����,�����&1-Qu��@���;�'MTy�g㗻��:�����/�k��qo� �p~�,��N�ҕ0�G�s��q����ˣa ����
�c���}���٦6��p��Ԫ춪�]k4b�"������sR+�0��c7�������}rX:��p�.ۓ�T�w����+����ml�3�CyRW��wZ{d�E���z�����RUUU7����N������j�5��ku��u����	���)|eR;�6��f�s�˅eS6���f�����
D��+`�+2�l6��-4�J˟
��fc���H�¿�i&��߳!�db���+�=Ey#����Ua`clO>O�.�)��M4+�X�*����`v�����E*�.;�����;�ئ^(���l��������5�pE����)I��pU�;n������lpne��%*�sxW�u|`�D��xh}0J��Q?~�y4"�a�m��<��e=��j31��?j��U���_�6�0C �o���~:������-�>Xai�h?� ���*�j���b:/ܻ����~]~AA���������08��Ԛ�w�ט7�1�|��ND���	���o��s��m9?h�ݔ]8��d��F�Q��4l��ND��~V�~���x+�8�>/����
�Y]	��V�֍x���Ǚ�~��,g䊗��8sN�r��F�����$:Cs��n���N�G��S�����r羱	��H�WWW�=�	����)�f�k	���Lr^Ц%U_1�F'���s[q5��P���|�O�һ[�xP�a�C��Bȵ0_#��Ȍ$^qm��S����o?�p2 ۮ^�[};�կa2m<��y�hi:�x%[��2RX+�}�`�`������e�a��/#V�be�Gk�^�	</�]����Y9�ؾ��{��;���DWc��B��E�C?��R�L	&�h��H��t='���РsE�PHP���4�`��8f����7��������[g�};��.����Lك��C�4�E�x��Q']D��^���lN7f)b@6s�Z�@��܎�/.kJi$x[�/&GR�@$����߭�#<�%ݭi�t�E�R��@��@�dĊґ�;/Q�S�����!L~�c�l�8N�z9� :"�R�-�W���I�ȷ�("��[��BBq6�A�@G���j~����~Z���-E�]��79�o��_��c
�t,
��fV�8�>�4���9��o"?�:Z5�l�������{\��?�"c��Z�I��6�ZS���R�ڃ��5�!-��O��;��T�Q�f��P��M���ڳ�拶��^P7�$H#����z�_�X�6�!c�ea"�H��A�w2QW��G )G3l݇(	�Z�X	��|��V��=��d��q��XP���gk���r�΄(�Z��?b4*�_��$�֮��U����I��-�8�#���:��N��u�=��}\4F ׬�Ѽ� ���П|���g$������/�:Uc��%���-���e�v���5Z�lJk�X'8r����^��Z;!�����N����l���42���1AQ-4�ט�\���O����d�h,����+��D��\'�#�����n���(�Rcx0l~b�1�6:׻x�0�Z&p�t�>-I����{���:^�Ȱ��JD9��5]�D�Xo���ײ��Ƽ�:b5����I��{�ܦy	��T�����������V<ؼ��$���3��rW;��ɔ��̥���R���5w�4�hDz�gGCI|�m'��[[{�b�+��22�q��?����n�O>>�Q��3��G�;5$�z�ދ:��WyZ��8�lA{�M���ɏy�w�����-]/� 'h�/�[�o^����4F$ �^Gn��`�u#�ZkS���_��Ϩ=�Qjڞ��mGVh�f�]6?�kI�N5����l�E�M�����=ڏD~%G�H��3*�ݺӤ�"�I`��'k�����GݾM[kC$�]����??�#�����ǚ%�rR}��)2���i��۫'0�r���q�ޟv���#{<������C��FC�돣�d�;��|��7P���oV�X�f�A��#Y�ץ�rD�-L�?y�PT���7F����7���R��/�x*R՜[��O�0��g9HY������*������"�9)����T����כ���BI��ͨǄ���F�'vɿ���04�m���:h#F�d��"�O)$`b�MI1��*�/L�0l]�������w=����]��*R�A����e;����Va*�@�`n�!\��%S�l o���0~�'�\ �v�n���	M6��t�U1}�қ�7OR3�S�4�v3��?a�c�y;{~�B��j{�Wn��ã��s�{H�u���PAm�_���ٽ����8�Yrd�ng��ApwJ~���fsZidܲy�)��\�E�a��dl0�4R�tE,�4ƚ�0�x�E>�>��wK*)5�-���K1w}���EҚV�k���LK~rzo��,f�[��9�Vd�ћ�☆\��G;�?$Pj���hT����R�c�z�D��a�u|����M u��=�]����?�0 $U�h��N���~�%�[KU'���L^Q��% ����+�ϯ+`��pho֚��_��fG#L�luv�sc-P�+H�Σ���g��ϫ��	
�#��4aUKWD"O��ޛ<m��3�U��	��Af���2P���Ғ��E�~��Z ����hī�xω����=/3��6X�WO_ެ�� ��Q�8�e/�F�D8�=��c�J��N��TOꆞ''(�D}��R��"��r� ��w儜�F��Z���mRC��/��t�2��T@�`��˻e�9��@N^��K�.z:�V�Fj>�6w>5x8�S�k�Ba�t��G�2FD#��Za�>�L����s-qF�sa�?H�%K�wM�6�Y������	���.-t��>=�iR�C,f��wc���wt�UO��9M�t)LR̓m3����+l/S	�<6�s��)>������{�\���Aq�_�7EAS;ܱ���WL$ztC�?���ID�+��!�+�bHV��N!�LdIp��Ǭ1j T���#ԯ���6����_.g4[��4}#i�v�ߞ=�&%+t�Aώ�I	�2N����'�[����R+���;���h�X��;�[^5���Z	�M�mMM��P�Z������� ��9 ����������Q%���|}�ǀ�c?i����lNg:�ɳ*�~��0bc��lVE�l��l �B�[�'H+_5�'�.��B�����[7�kEH����K�}�t����؝��Ȥ Qc`~�7�E?��IYy�� �ֻ�5ZaCK�t��i�`�gv�N}kkk]Ss�N���{�Zu��N�*+^5f�Msh�g�|8����M�2��_=e!�;���ɸlv�7��_��v��M�(|�6k�X�2����n/*� #���eT:k�"�wp�p�'VM�6����0�J���۵�]%2/�&�^�:E6��E��T�#�]F�{�1fi�@:����>�vU9������jqϲZ�/���<������h�qq����n��%rM�j�۪ ������88-S���C�D��j���T@��sJ�7�O���,0҇��!����zP���rр�٤{��l�ھ�T;�T�!:��/�<J��&��i��-T�r*?~�W;RoN�Z۞^`�4fd�[�N#����1H��/�g�qթ�9Ȥ� �L�&ZP�\������#����5�:�o.�&��4�$�ioQT�X��B�¤��~=\2cgO.�*^�X��I!����S������+��ܹ�y� �ޟ/4b�n(�$š�?рiL#�ؤ���RG� pQ�8���ı/"��KG76���"l �	z�g��Эq�UV��?dX3�%��
>�>�,_c�)�}�
t����D�4)2��7zN��X���?�N&��s.!�����'���
bx'oH��6,��N��G8�(�&)��q�)~4r���qO:j�PB�i�&�L_���?���. ��d5+���t�Z���o�Qٵ�����/;��ݴoo�GG7,I��L@K�S)�֫���r�>�����������V7�\�[1R�c�z�A<mS�k��~��א8��,�,P-�7p�T|Ƕ5W]k)������PΣ�ū���\)��`��Q��=(�cNZR���p����p��! ���~L2��/��M�������Z����QjUgV�@��ٟ��"q�U�U�^�ۮ�m����B�f���|��=�-����	�M}	�.x1�{O9��L����y>ZB�R��Ô��F'�B{�
Z�v�NP�s�t������_���.ȩ�� P��#>���_�]����>��ʿ�q����/Oy@��x�4��="��_	BK5p��v#��,���h��4������=�F��S�Aۿ�p�*,�������'��p��#�H%AowS>�r5B��L������z�W����gg�e 
��s{���r��Kk�����HV՞K:>�Iz\�������wYY�c.��G�������]��)&���T�9N8!��/R?�H��17tK�+�1�5�.�Oc�E�Yr-�',��Ts�����C`���nl��C�~]Sk&p��c?�Z:Dp���U!��ۇ�8H9��x�c����%i7F��d�<�ڹ�Y|�0迎D7hu���,},�@�_����%�!l(A,zz�(Tm�b ��5@��Y2�bx��4�"fMi����)�,B������`�|��ޞ���(��� z�8m�F�{̭��vOi;z�����Z�.:�z!��R#����o�������JO�s-�n0�Թ�C��}�y��9!�g8�+������dwVmuꯜ�q��jsq�qs����X2�{8@�5z��Ub8.J�!1W�B��"z=-R"+}�]Г�V���q��A QVv��ڪM�@
VH6��,*�KO�8䴳(�^
��XU�r`}4��ϫK�__��Ъ�ӿJ�:���^�p���:�
�?g.
�}��þ�~�)�_�	�V�QٰcG V�*� ���T�2�F$,�>H�h�Ӏ`v W�]��l�]�
��m@r��m��hzJm��#\�����S<g��/z��[��H������ɺ�LE_J����|�g��ƌ�A7�ھ��V�g�Nו��� �ˬ�t�WЦm�3l&�)]�h���t�3�D+}���%�gM�f�]q���j?�~�ދȣ�cX��8��w�n�PfPt�|��%�sy�:�N	����"ܻ�L�S�#pԜ��އ5�,�O�O� FH����T�[��
����	P��I����$��T���x@嚕����ӧ���z�'�Z�&��~�z0a��t@�9[�%G��Q���r���b!��D�-[Q`���'4~ld�S}_��L`��<�����[��a�W�Ŧ��Οģ/ځNh��Z�p(X|1��8s�Zx �-�A�x�ʝ1o�t�ʿ[��\C�ҩ�\� r�K�hPuu�������eĩFDB��R	N����,� �\�}O@���������"�F����O��.E3��pG��)��s��Ȅ��P��Or�\�3ۀ�g	d�[�Ag���U�hE�����R|I>�~ŵ	�߸��ٲ��7n�5���fd��X���O���D{���5\�G �klBp��Mv ���r��? ��C��(�J����)d����BP)�U�y�C 7F(�����g(ݨBN��=�ѹK{�5�7S�g6�_7��~�rp�J�f� ATj��
%7,IK����Veh�r�a��<�p����d{�d{���/�M��c��m�~ ; tE�tp�돣N[�p�u���a,ep��	��t~Z|������I1�s��������\d,�N�HZ��W6묆d&r�HhѤX�|T�/��vPk'lS�?���	l�K�"�X$P�c�%RtM�&��c�W�8�ٔA��$Z�Y%����4��	[^�]L����Ԇ��џ�vw_sQ�����y'{���^�.fp�Ŕ�"6�}�liX���j���v�+����8H]͂Y��>����ĢTiJ��	���g)6)}�B+�߿ �04-^ı,BO#I�PPP��ugUh����r�t�y�/-���h���l�ٸ������3�3ᵅ�a�d۷��h�;:�2Z}��aq<sXq��귌�?��Je�`���M�vI�B%�M./;L�mM��7`3������5~������f�͚0�g="��4ʧ\Dr[��Y�[��O�ݹ�˴�P;����_��>��RO�ٔ�bX�� �*�=��p��p|��'�k�'P���̾{ �6����ݻw�0��U�[;��{�㘋~وA܆����m���ǽl.cT�c�@��.ES��9wk��g�2K�d���J��Q�z��!,jR�_GA��;��;UJ
 
��ƈR.]��?�g��/S���A��C�#Nd�Olx v���a�h$�����_�H«(*���Ř�K���D�-L��{�b�[>D�ӝN��a=��F"���^&$���C,0�կ�����[���/��V5��T_o�����FĿ�8�� &�@��bPw[�������i��eh�A�4�N���T������}[�tS��Ѩ��x�Ъ�e!�<rؒ����E��'3����ǧ<�%�/>�p��]iz��7M�1~v{r΢���И��Ŕ\�����lU�����B#9fn���s+������tz?(���p��`�3�n^�]�Oүç��=L��?�خ!(`�=\j�I����A��)�ޚA !�X�eZȾt��1aͰb�S�ܠ�3�zI(�ԓ�仢���:5h���J�$�(H9G����HX�g�434�A�,lk�*�5|?�"��<ʬQP�y{���$��45���3Yvf X2����Z]B>��~l}��p�	J��-Κ�'P@
B$�rn�y���Y��~[;�����~���y�̃׬��rJ"gb��D�9+����KY�_(��V��ڔ�.R].�.�Z!8���ݘ��`C�S�z)���>��ٽ�%?��jn8AD���״���-]�ZX���~. *m�NS*��,za�O.��&h���W ̣������R˚�L�u��oA�Nc�� �K�M�/�O����64yL���n�.[�D2ڬ�͈���S�j� ��y<w���)��}�.������=҄$D�Rd�ԉ"߼L6����c���|!��\�費A�4�rڎ-�Ct,�ct�y �k���R!cT�|��蟶��E���XR$��@R
�#έw�.���E\#���4gbv*.z�Rc�T7홏��I�د#nt�����?h�=�,b3NN�l����c	6�׼M>������Q�	.���SK��x	�a<B�E.�Z�]s�Z���߈��� 1��֐�D�=S������T����V2Zf����H[���ZE��\�"ԕ�F\{��}�E�-���е�_o�����N������|�����B�T�����Z��KS���<�?�3���%K�V�A���+z�Ϥ�q.Q��':��?�ُ�=�׿��84>ZA�.&�
��Lw�!\=�3�=��'Xc�$AЙ�%����1�ָ����^���7.w�d���C�),��I.qʐ����{߯�c ��p��ҝ dj|�a�� ��B����Ʒ#��~��}gy�oqg7�C�ڌa�m͡�ÁB^y����dv�;��i4�5��]�\~!��Q����<p]žEc��>���P���c৞���4�8��̸�-����L2����f�;t+󉦔��F��l�dK����,�ݡ�c�pg�E�iR���#T�/��ۑ���fQ�)�߈g�����^6�3����!�bE~�&��ş��X�ؼOkג?�����73>�����
Z���u��{�旆!�������oP�ܦ�j��0���|)l��S'`S�P��?�S_s�p��J���9����d[�T��,�Y�Е�{�QW����<�G\��,4�i8l�A��͢��Tm4�C��3�P�$���g�CE28}��З}�tZ,�L_%�~�Qټ��]�F�cv"T_�:
5�օ٬0j��S��m( ���1���61���2�)�৮@>|�	X�[51��;XSwy�QG��\a�u�?ſà���Gg��& �f�Z�% �Sg	�`B������9Ȇ�Ш�X���7��x�d�	�n���!��o&�P.��.�ڮ���e��
��K���G�	�~V��}2*c�UC|Z��Y�����B��$��F�5 ����7x�jEct��݀�l�U$]��{���"]5�~���B]#4��acN:V��OZ֊L���ts�Fi����5���	z8�N���4��2RLD����1�u��~�����{��f���,;w������Y.��aX���bE��������F+��n]�/5�����>y�[G�z�J��f�!6/|5iv���h��Ȇhሃ�;4�#�}�������������Fb��%;��DI9��,��ڧ��v��]�,�z�)s�97 2����DLQ�dKl�U��9!HoI��ܓ��J�.����E��ܜ�[���T��{�E9�c�����W��k&�/�CշEA���=�%W����_.I�s%��~�7 \�:x\�|d�U���W����c�ey����'K�._����B���/b�����E�^O�F���"ԗ�"�� ������>��h��
]. ��ؕX�H�9�E~)z�ցb��0��&�LŹ����_2����\y*������W��������JQ��dpvr��S$�,I!���r��띾�h�&`D���&�;�i�J3����F2jcû;��Žėc	�>g�c�ZZ9��O�Ζ���5Ł(���T�|����`B�`*9�D��7
h�������1�/I�e��4(�$b2�6�k�]���:�y��@wN���B�f�ϒ�>�(a���>W�=��x����R�A�{8�3�����/�C~�4:
�8�^ӈ���}��:c3����>�"�-��ZhKЉ8+r=fj3b C3}�_����b��c�ae�Q'w�2�BefJGcP�c�m��Pz�q.t��`�%׼c_;��?�]���q���{"�wHE3�VO~(�|3�~�j����.���g�x�*��*,G7���3��q	/�Z�:� �uh9fA�Yb����@*S>F���>:<�i�X�I�-���W�����/��>׸Ys�S��7�7Ug@����h�SrJ���袅����!���>�&��M(�7>����l�^�H3z��sj��g������;��,4_p�DW'g��;Vfl�t��|_[.%�m?/d�?���8J7Tor=8@:�2(~�(�R�W� u(	���W	�Ǯ����`n\<p��B�
�-��~[㪙��s�`���]o��$7��O�v�G�<;h0��^���S�_)1���>�u����&�+��e,�R4�:�Eȓ��W
��O��$���̠,D$x|3~�~+�/ ���ac��$R.�:�
p�7�ǲn*�:�����i4Zjb��k��rJ�:�>o��R�U��hdl"�P� h= 5�k_�f��A�6TJ��	��R:4�s��ZvO���M����K��5��O��3`�X�y�y��	��I9"^�E�Կ��x�g��@,(L:��,*�n��s�$���O��$ʓ/��
���2O���=S=�BmBr�a�!Q�?�n	�٨h���������<(�x�~G��0)a���bXu1��p���"g���R '��������E#����=���**aE��O�����~6ό���׀�u&�=�и�<`�գ1����_;�)Bc�}���Э�~W�)I�O�a�,5*�*,1�1��a���_��'�I!N�Ms�f���ޙO�;v�-�p�?SL � t���U��H����\�e'O��%�H�E7��#E��H#�+�>��ܿ�cH�j4��cȴ1(�
�°�t�)z��;P@5=�H�?0y�$b>�)&�S 29��`t��`K�T�bqhss�}���F����|{N��p��r��L����L��f�:;��sB���u�����,�E����+���z,5Z�m�Q7��\��}�e�B&�0'���p��-N&�(�l����?&��āl<Q���5��c����i��w*��iSrf�wMxI��UN���W>�s��� .�"
O�d8w��er+����rJ�R)�����1¶I>�D�8�<X���:�_5IIո@����1sS|I;6�RDq�: )�,�3m�p9'x14�#���ƑOY'��!�9t�5z��5"F�!�����;����c�9M�wt�����8F��;Y6~����J9� �BY7t�+����lY�m^8�p�,��E��X�d����x�u[4�7�8�
h���"���� �{��w,,�;���r#�S61$*c��IP�

��И��q%��Q�$���`__��X��a
�M�ad&$��ᑃUd4�c��9��A���{I�;�����ѐ��$+��@������v�.����&?đ0�@�e= kj_m�����xX"t��$���bݑ^�"��������@�+%�Z�/�?mѨ�֝�&;u⡦�͔�{�=9CE ��
�Ñ�K�@�@ɻn��X��R�t4��L�zG`�ba��D�S��w!���^vݤcoBW�(3tX������Rʬ���Î�^���JGޞ<Q��s��e�9��$1I���PRTU�{d�����7�[�˷�y?Փ�|�I�XF�޹j\m!H1x_8R����&��N4��U�"`�>%�Et4X&��G����{�w[���}z�
k{]�[�{�0^/��u�[-L~B�:1�;m�\�IkO��^��@s�"�p=�*@u��'��M�˙F���C��d\�]L7	qp�}|�{��1/��'�G�CtF�ߪ�L-w�}���l��%���^J^�ey��z,N\\��|N�i�WT��Β;����B�T�e���k
���!"�P	r��vbV�yu�_�]h�%��K�m�f�����Lx\xZZR}m63`|�J-9�r�N����l�{^�9:��U����i©�'�<�c��"i�<�,`�oѦ��ﲗ�y���Nw�Hɾ�9:��}ΊH��p�H6&��54ۦ�_9"����+����t�l�x�ĭ9pp�J{�}�p^�{���J_2������/P÷�
������ ���5�!s�:!��l��'�L6s8�*=bʬh(��ur)��$O/�H[z���C�>X+�Q��gX?�E�z�^櫳���`:�38�(�r ���T4����?�P4���3a�!�K�e_��m��2ƅ\Q`{����wq#�o�������T���w���WS��(�h�QqoT�@K(1J ��&Fp���`8I[�I;i�8
L�K��~ʀj��ݻ�\WJ|�V�/����}����K� �"oh�SH����_%�Ţ�B�v����w��7��c��6�ׯ�c�F��۝"01�b���"���B���Ξ������.txoj\3��ãz�O�hB���qYG���{��(��d__�$�����ih�F�l60���U�8׸�F�!/N�PM�����G����@�o�2�<	=ᾙt�6|�8G��z8�v5&���(�ިq�⥠���N߹�&�&J����:;!����Q[7�)���(��y��

&������A��]�3@W�Og0����
���J�-$v�B3~b�2b�|��i�N����,j��ǩ�����w��0����&��L^$;��
ੑr��D���dQ�S�+ާzUu��S^�?��]�@?�Ky��*���4H�L�8�	f8[jp�B�/~������.>���b����|"���q�.�5{������^�'��	���m`��jz=���-�x�*z���۟gd?q,��#�X��(|$�p0U?��-�g���E{����er1h�?%*�H�?B�-�GS����]Q�/_�GU܆nA*����;W���Ls���!$���C9ڱ_������"O�U�H�& �?�=�_
���\�zd�A�)��㗝	��7Oz�:��׍��3�vjJ�w�z���ئ?F��kl504�e��{�W�sK%AӉ�F�ŝ��w���ûζ.�����D6[�!C)�^�1"S���L�#�`���hm�荛�Z
1bv38��B��>n�}�(q�TQaoc�+t'<��ߣy������/����:텒�Tg)h޽�p�� w�=�K��7ۗk8e�@J�"�$,�&���=�u�{�tc�7fzG?���ֱ��j٠�w���j{�Y�kO����%8*w����<GR�n��hc�n���T�/�W�^U�A�h·3�*T �TK����W?��J5���D��� _�E�{�'8v����	��&���dI9:'��As���^���(�Sm��]q	H�#�]����!�
��_���ip�B���ÝUA�v��,��~$��aa������9����_8����/ۧ�������_?�o:�|���ၽ��2?8�C����	�}x�i:[��y���0;�$��'���GSߥ�Ε�����/�w����<C)�g�*Vy�����c�gy��ˢ��dgUSc9� dB�2�۫��R�ˀ?��(E����m�V�st�uZڝ�P4������_X�N��(z�MY�sM� ]�,����$���$�����:{;�UC؞�s��e�Q)$��.�8K�7
��=47Ϡ�憊t��|��E�=?�����KZ*�=	�ޠ�s�:��l1���R����bj��T�>��C����ZJ!����]o���(��"�_�|B�ك�����G!�+f@T9�l����A��� C"��N@���9x� ����l,�����J�0��������$������w������H�{l�,�e%�L꽯8LR__ߨʈ�̚\a`9�Z���c<DBkk~����=Ѓ��s�%�=��=��M�U$�W��/�^���-��2�v��u�)�)��?�Ru^"�Ǭ'��#[�:;M]�Z��kh��������7������Z9��ٗ�De����N�'x�*��^�~a�����f~|V�+��řw]������Sg�ST�vZͬA�&әq�*�%��T�vxx�a�֏~���D���v�S�`�ꂆ=��6���_?�����W����H�h�Ba�����!���4{"ۊ�i�4~J��+en2��Ěf͋>�S3�� �j����iF�	�hP�H��-j�oZ2���1\#���N�M��l�]X���$̘���u��7����&o��]��n�^f\(~q��֘?�����ؚ��������)�UiQJ2Qq{O�0'C_�X�NO8j��1����A!
O0��A[Z�\Z͔`V�>Kj�/��(�E��bȖ����MD�S���K�Ey���b���VE~v1q���歳`�*w�oZ��Y��߼m�Pv�P"_�x�n/j�=N+�5����ϟ༸q�Gc��pt�z^�lR�,:99i����tdk'l?AA���Q{��wТ� �F�.��>t��^Ԅ0#��h�I�`���r��7F2���G����[MM\����#Y�d���|p�4t:�5P[8%�'�P&U�vC[�B�N�)&o|��&&&B�@��GB�<��Y��;�iM'$��,bo���MXCa�t�!X���0
WuA��s|L�G��Ci���^8v���Q����4���5�i�`/2���	<��SE;t�C��D�@����4�U=l��z��Аe!)Ŕ�"C���P��@��s~]M8Z��qw���o$���0a��go�׏#�s~��N$��"N�b�uH�x��CӦ�/�F�j�У-EEE���<�U��ΉY�R��;��c�����
߉���_OXoŻ��(~j��5#x���;CΜ��;¢P�9ă�2����_P��X]]���}�뇡V�o���D܍ T��|�����ih��0-��
�6ι@7��5�!Q�#5�~x���w�l��y�꟏����ە����(__��������j�%q�y,4��nTO(Yh��o���/�㷭���f��{�>ڛ*}��l^↝�h1�|���O�K_��]#))R�Ss�����}7O��,�j�/[/6p�P1;w�s�1⛶Q;��lS6޵0�?�}o`p�>�F�����N��88^>�-�[Oh��+)�k,��MD�ׇ�I�S
`�,�T��nJ��+��|yMM��DJ��j����� J������ǀ��� �O7Wr��!�8�69C�?ws��~�����&�Uό����3�/�Mĕ �i2�m�p�z��2�3�A�J�F
+�B��D)�ǿgS�e!���$�L���Ϧ�{���R�d�7p�Q��LM1M�]�:���k��#����[�܉��V��K/(�ry��`V�F�l����ki�Έ� և�D�zf��!��GM���}�!��'/��K�<�˚�A=�q�i��ё�H�:���h�14�7?m�,2/�_Z"W8���X4Λ��Ѥ�ݺ,�;�u���$��=U�L���N����7�I���V���o��af�,*H��m��q�\��ntM)c��#˕�L���w�gk�J9"�p���g�m���$Hީ�y6�  e��W^_��ӆ���*R/o�7���LS�J队���T��_�A���*�|�>e��yۗ�cT�X�
�f�o]�N��N>V֮��˗G��Iզр������(u�2*i�w�|
�R��s���P2
�f���̑Y�8��KY֛�
;}ӫ���_u%r�H#v7�-|��1���V�1��T���3�&S����-��~����[4o�zz�n�rwwO�����ո0�Omqx����~�Z;��:�Ȃϻ�ƅ�;�����I���[���5�1�R{<�9���~¬�0,<q�{� ���jd��W"F��t�2�z���^���7�*AF�k��zt赙	5I�� 
�M��'-,|h���,B�\iԱ��nuR#�͂Ỵ�-�#��8
Mu�'?�:kk?Yr���P>;�I��U��� ���a��Io>G�ڙW�5��՜�6� �N�k�h,��W�m������	xإ�2���7%��D�+a�"Qd/�;�x�3��O�c�7�O�GAՐWP��"���ق_�/�^�)�g^��!�OL4ϯ�Ȟ8��%ti�"�t�c�f��&mn�Es{�b� bK<S=� IG��jהOm֗�KZS�20���<{�:�h��(R�~��1�N.f<u=��b���)�W���_mFpݩk{��B���ua�~Gm?��n��K�t��A�I�������림j��&8�"8R�;�[�n_�L*ICS�%��~?<|������0���6���R:���qN�Hd��`�� �}�y�Gt7������D,5Y�8(�2�_[�B�W3�8���}8��|��#h�Y g����`d:KA���p��N˦��0�ε�~�6��jm1ֲ)�[k.�%Ś!�fJ��3c���tC�FFF��m� ���B�N��Rf?rd��TG����)�����M�D�H�.�s����A�qXx�Z"��ن��Q�w�ɐ~4�`�G�n�ӑ��1�~�<��Z9�|��37B���b@(;�Y��x��;������mL&��k]U��\�媦�F��s�20�����g-N�x����6�;�p��`���D���D�n������L�h6[7�Ά3�l��q>8�g�c*��J��ۚw�$>)���?������}�"�h�O��0�ą�
��N�cy�L�ΕH�� ���?@+K�|c�|�2<A���Z�G�тn�ZKu|�ds��E$�U�a��8]C+�2���p�����5���������E�sqX���7��!5��g%�{>|�.���#<��A��*-vzEO%~n|��w��i%��&���T�:�'_�A#5
Ŷ�{�����m�[.���������{�y A;�׃4�V��`�0�C�m-u��z1&rf*v�|k4?�zGcp��]����@�4��zg�\�������6�{DN�v,I�^Ki�aV�G�Ld������S^�� 5Qvt�o���+4%}=f�K�g�������7�൪p{v�%�瞱Ǭq�8�&���\o�UR����~���QƗe�[f�����RQJۺ	��S�a�JŏVIۯo4�$�)[vg����6?�Z�s�y�޿}L�!k:����o,]Vg�����<���q��ӬϰDlm~�m�J�Xm)��Q"���+w��9x�Q2��xskk/�壍huv�t0X��R�[
�>����-�a7�Q��ϴ#�h�� �k|�M�WSS�WǽX���'%���_&�.^��+���kk���>���g�d�~�鹸�FKٔ{�8�[�L��l{���47����5�yB���V�ꟗ���D�;�$t���/n7�+����9xvѩl��(�����2+��%L�џ�J�K�A�*�ڤ�_��6���=����[O�b�&��ws�m���"��M�� ��#��n	�d�:2~fN]�фh	��P���p!����j\B)���!��B���9]������O�ɚ-o����_go�Ā�	H�J�P�>I�/�q4�Q���!����Ё���ul�FU)jس��q~#�[��]�'���<mV|a��/����eW4z5���(�n٧V��T��ߴ��^�i�/�^�EG]��G���޹N�~�b�K���M�5��n�o ��7�_Mp�E$�6�c!ͅ][�n���JW��^�P�B.@9���e\� �A�6��Z�K�x���b�MsGqx�:���k����ƒ��h��
n_��`���qr�PwL�m��R�Cy
�tJS�"�ym7?r{d�t�ٻ.-@�:�����������,�7B���$��9�u����X�X�Jyn,�ߚ�1|������5#N������5KLϥ�e'�mb�t��^��Sm�۰�[���[���]�����U/�BSc<*߄��T����om�s��\dd��D�����R��=m��#�q�Z�����n+�����e�L�_�Q����dk�b��+�-����H��X�ۙ2�����ȭ�yU%����t��Qz��*��],� ?ou���^���Bn]��1h9��T��D����I׆��wC�Dlv������s��sن/J��0�fz�I�=��Ԫ��G���(TH1��)Zh#kt�R�`�4� qxtѩ���#��2��=�E<���s� `tE�>	���fӞ�y��'�΄\z�&��Z~t�+�ўX�|Q�/��l��D_Vh��X�S�i<;��l���l]��97?P���r:�C�_j@�Ve��ȅ��o��ثu���R�ᯚ6~�6=�җޫT�U��af8�����~_!.n� ѤN�S���w�8�y�m=� �rۮ�YS��:W� ��-��F�$��D�]��7N"n������`��M,�Y6Wۻ�Ԣ���sEI3����oztˆ��ԕ@����g��6��h�>�n\BiZ@}|���
����vvBs��w�#�`B�v� 4-���7%Ƣ`�����{,��V�{��rW��}2<@$o����:Ԁ�����"X���z���\�CYF�+TI:�Դ��O�����G�M�2��u8�v�|j�H��!���?�d��}�O0Fl����=:�G�}�C�){���ѐa�,MJ�Q����2�v��P=����R�����ϗ"}�L������!4��`oME�S�a�[��y*��G긮}.Fh���^桇��&���W�աz:;���K|9���#��1�k����Ҥl�>K���=����j'n���|q�/�bX�ܛ�l�QQ�۷/������tR����1�+��ܪ"��r󡎀��|�����*��٧��	�I�k=�V:��!���]p�kN a��$<�-:��r��#R(e-�gI�
�AIiiO��qO��"�:���x�!߸�ܱmm�'�˔F0�yw+(����~fy������[kZ���n�5�_:��]<<�i���哪L��.�v���\�����[*&Ĕ[���{g�An��Tp?A��W4�g�Ζ0r̋\J\B�����|���7���7����_n���O^�Z��\�L�.J
3��N���aI�;!0in�Va���{��&�����K(�0gd4��|�h:��k�K@�O�d�m��J���h����ʎ�3�l��ZӃ��WV��P5��xئ@ڙ��*v\��gN�g��1 x&�F��'��aE�Vyj�{���>5%�3�vٻ����{`�-N�)d���}꣬m]��P�i�V��<p;�񿴟|������b��usrz�3'�զZ�xH���&�ێ����V����H�����V6�w��x���S��S{j�?�ȼ�_�}Ɣ{��a��yf�M:d)v-:ￛx�Q���*Pp#J��������Q!��V���w��9O�4ϖ���1�>D�S/�����]�������H�%�>]���b��J�[Y�ۥ�sN1�����ݨ�/&0L�sy����/�^�	����*����֪}t�5�]㯉��ޱ��Ah\���ݶf+�3'�bemYEr�� ci�^tdѕ7l0D;o��vi��w��&�T��t!�p5k�K$�د���4ߕ�Ȇ��x�/*���/�����!sDg���~|���ƍ�/f�	a��^j��SiD�J��p+�^�		W��(��Pk��Ly���+[`#{6I���%U�r���R�/o�%vQ��Z/lv1��Q�`�Qv�J�hsrNj�Ϟ2�ц����y�W�c�և2,�K�;F+nʔ{�2J

��3�Hc	�R��$G�BF�n��ϓ	�AO?��.��N\ӶT�y"z?a�м���ߊo�@������~m��a&�b�����[+t�:����@���8�3�����@�#����{8��n�TJ��XbxR���?!�+nIl��1�����wG5�@��uTT��4P_��Q��r~�	�qq[����F4��Q\��ص���ke�������Ҳ!��d�6�:���1kݶu�X1�1����m�v�X��(Q��\U�p���������+Q3���y[�[V�>^HLז�.͛���֚�r�<E�F���i�=v�B|�5��k"���w�����L���Y�ؒ�z��3�{ ^��.��k(S�9O����6�S�([��,�`�]��wN�%����H>�?����|�r����6�L�R4��_h�Ҁ�DG����ǖ���C/�B��j���!���󹓓�r��/&���g�V��e@Ơ\۝�߭�{��Q���=�� �
fo�6��VL�)����K
�WU�-�d���Z��z짶���A'�-���im�#N�h��ݛl�49�`[�����0��=i2
���8z�pk����"�U%�#�d��������5��b�3�@9�V���Bm���N�e���Ύ�'ۣ�1-��=�����l��	�5�;�$5��=���c\�BSH;2�v�1&D-sz�:!Y�]�m�+)ϡ��O���ʚ�w�R����'S�U���~�sh#oߠ6�;7`����ߗ2ͤ<^8����t��H�lL��M�=�����+g���({{�ܱ�k}��3��!ʹ�΁k5�~a4}��!��₭�	d�^�_��:ў�n�$���!j�Y��#��8W��/y=��HKK;��%R�KC�]s��R��C�\�.��9�ݢ���te|/��J���=���8[ xff���X1
7_X�EL:kQ�]#$xS`�l[j�M������*べ��u�������ܱ����;&���lgV���**'C�S�_�O{~�@}eP�3QU]}6�]��v�����ѽ�I��]Z�<�'ݨ<@�`tD��KJ],�̩EO��mʕ_H�D��1U��?NG�hM]�ϱ��\�iK�Z�k��ы�ł�'�W7Co���:�`O�Ng0vvu���Zym��^�;;9U:�d�.V}�H��������d�%Q�����/�ɚX/��Y��8�W{�@�s]�K��5�8��!z���r!]	^w򍍤�Wv����O�a�������<�$�8\�=66�r�Ն�iwW`�fi��v�^�/�����iY�Js�X[g�8�������S����j�Vs�������������h(�^�Q@g/oР���e��� }=��X���й�a=���p-K�����l�z�F)��T�4?ĲdX��O��<k�r�J��>�7����o�=���0���P������J��ö�]j��?C�lM�̩�6��u�PҚR딗��d�n�91���
��eϮ���t-��?R3�S��4����G�YTm8c�N�[�)J�ν������#U�uuuМ|�guqE����b$�-	4����9�jJ2V��Crn���f4+6��>��GP`jjj��õU��?�_�h�>��㙪��k�F���p9�:�����_�ɘ���P�Q�Z��yP���N�S�hjc�ۋM^��t����맇��ˋ�/�,��c��y�,���s6��lv�9����tS�����
`e�]��(]�P����QQlH��� �U/}6ܘ�h��R�9mĘ�d��f�$���4�[i_�]_��)�tw��)��������/x%�߅��T*_O�b�V���}J�س�j@9��1�����#�2��μ��sԎ�l��4��TR �~j5hju�d���|��O4�\`�4���W����0P333#��J���eftv꽯7a�C�&4������@�QhR�6Bj2�~R�i%.&����m�p��N[��[���.���u���� p��sSRO��	`Z]�������tG�?i�����>H&zTKxn���p6(!o�_u��d���:��3���5~ȕ���P��d�i �2d�k8�~Q\]/;���iy��D��_]]��g����� ��ۗ������f���<q8��?�j^'{wgN}}#T���	4s�sV_�\�{Rô$�4Q��{���~�q=�mJ(QU��-���7>�p�a�jUԅ�Zf9=j\؟^ϻ�sK�Q�"f�\k�[���_����ƍV�L������J]G.q(ΰc�^��b�@��D�|�׹\�ܭlI剉�@!��a���gΜ��033�sT�*�� ~/�2�ATWww��pCn.�����yc�����������Y:��glH ��+*)�?{v���,�R,���L&���H�3�b�^l����zzzofX-X�̡�4��dB��v<3���(�>=5777��i��-X��ǂ�%��� �0�2c0|�~Sߓ�t����O�r����ϓ/�Fd��K�`�c��s���z@B?��z����($�A��x#G��nF�:d.� �b��J����V<��Hv&����lgCj�i`���Q˻�űB�m�#Ma��r�TjKu�\�ˍ^��s�$+�Z�A�	��ŕ�/,��1�*��xM9M��G�d��d�A�W,�5�M*��þt������8�\�З'�ي�;׶�|�������(��� tv��ܼ�����&-��?��?5��LWW��/eۮ��/�er�G�:��:- %��y/�<Ew?��j�R����ِWZZ����K��}����ǳGmI�VZ[[�Ԋ~����^=�?��Q'���={����q��{��@����su�N�]����h�$������{N�-��'R����[��ͱ'��q��<Q����Q�B���A��%����n%u��z����͹�v���\~�&ό��o���j���gS`)-��"��	�����9b>�
�OX/�Rh�UBq���3}��J'�����0���'�*  ����^��b/rC���;��/n�L��S�cf`=��Ҍ�-�M�nħ֦�~�c���O��Q }�����H����e(��q	�x��E"��R�|�
᭫���:���߫s�\���y9������(�]��*�S�+=�9�N��瀱��������a�I��{�6~�Ħ�-��Qi���� ��&8���db���p�唕�?~� =ǹ�����Z+/$�O}ȳOT�� yDvnI�Q�X���Yu
f�]���V�5^A5@�u�Β��-3Ù'��@� q�T��g";;� `���v��b��Uy�����.�H,7�ua�[�4��ұ�þ�$��ϋ�a`��P����j�q���[
=#�L��3YJ5Ⱦ(����o���{�x���}�Q��;�Z�K������/ġV�ΥБ���phMΞ�q4�ąTbk����ƛZ�M�� p� ���wOO�l|��ZM�B��!�%ڷ�=�Ll~���5 ��� ��3h߸�֗�h<� ����鹨Cj�t}/zf���̀t4#~���P�!UB�X��6	��K����=���&��,�v���-;�e	�r
��uF�e����`�|���o�O�����P�9�6�W�RI��Q_�m���C�:
�������2ٶ��Z�U��S��\SR��#<L�EJ��y�yM�蟹�}��M�{�4i�2�>�|V4��].�B�y˜[e����"t�q�_W|ȅ!u�U���8��Lmm%55)�_���������Q�D^ޟK��T!���8Y5�����@6����
=���g'�{W57��5U��vil|{��-����/~ �&��⁢Ǐ_��>��T=�����Z"����5��#��>���o�1�J�[Q���|7n��>N�_�	�f�]�Zm��� .�'�$`����!X�Q ���n��5���X�t�z4T?"�T���,��2$��K@g^������h
���X ���r����a�aLH�e��АÓ��p�r�8�rnccc�u$Z9��$�Ӕu؄7� vf``xY+����a��[?��ɇ�V��� `�$a��ڀ�{({�b�����UFɔ����І��Ng����������[)�p;"����ҷkg���|�slM���-�!�a]e��>>�@!��mU�^���0�+�Qs h`����X�J<��c�0�}�]^.@���tfSvi��j���/�Å�[7u�;�GB�WM^@ɿ��Z)8<�7�r�5��8�����,s5��ҷ��,���M�@����;�œt�:���Ҳ�����pN�tT&�}�~mt�(X?[������j�¤k��M���#����+�^~�F\i�]eGj���ߙ�,j�8�|ȍ �իW������d_(q��xω�@���F�~]�^L��������{MK���><-�&�4��4��K�苖٢QQ8���%�cOJ0C��g�12r58����텇��,�pa�o#��絛lJ"�n�>�tF� ����JS>��O�@�2Ny#=�׮#�!�y2eM~�(�,*(�x�?�uU+�=\�������Fȥ;8�{�ahO�'��痖,""�O��Q���'�T �E����h@�^����p5��H&�TV�q�r���\MG�y4w��V�R[�=�b��a�I����qC�U������lH���}�|!�뒂Z�t�6�Ԑ�U�_̢cZ� �����S;�n��.����j�CVҚ'"̊�1RHT�b��죄����Zs��س�I:�R�%U�%�E��섄���)p�;v���g�H��������2��Ѵ�Q��� ߛHUn����@|��(��6�C�Er�^/_uQ`C�7��Y&0p�_��p���P��*dR���u���!>�^������	��k�,�^yM0QΦ��RCbЩۉ:?��6g�Nܱ��򍃜��_�Ϭ���[�93lcE���%^����	�܊�S�ڗ���Ԓ��#-�dX.�j��ȡ8״M�Pj�{��� 9����YYZ:��t����5m���7�&B�B���ˠګ���y�ܚ���*~1�O���j�`*�F��Onz�,sZ
�%A9V�6�,�E�+~��#`�r�6a){�������^,���
(K���f�~���. \���,��ڼUUgۚW8O�z�?���X$�c�B7?~� >��e�5Q�驏yB��Df��I�<�KĎC^��.n�C[�U�xC���g��l�`϶����a��{k@t�	Fxxd��_��h���u�
v���rHc(��z��̣���4����Vm��E�մR�B�02�s
֣�߰��C�lWn�\�S���#H��s�{�>�M6(�B Y8�;�y�>e#�>}��l�(�v��	`�g�%1�y�Kp�T����<Û#'���A���a�!�7~M���o�zj`mt������+t�����X/̞�x��%_Dkjqkj=�y�IJ�Λ�+ŭ���u^�5Slp��mwww�����{�](��G�wG5�m_QP�*
*M�WA�tD)�"�z��Wi��@��Co�ti�w�Z���x�{���;#��:��{���<g��.�H��7���Ձ�'�㇛^G&v�G�z��mV�u���X�A�C>sraX$����f��"*Ɍ/@N�8+����3i�Z}� w�j����g�m����$��;�Ȋ�i�	���˂��l��:�y����0S5��ͅ�Ψx�D��-99y ���M/.5
&H+mDx���y �@^?J � H�p��٩��1�tM5�9�����>�/W\�0���t�ޣ���vu j����>��8$K���A�%�DtC=�&�>Ѡ�?ծ?d=�o��W<_	�P�5!� /����̄�����Q�A� ��ҶṺ�����k�U%L�=$�g1��؏>ܨu���M�}��@�y��
Xxtm#�s=�H�!���&~�r1��=mξ�)S�ֺ��H��a����/�dn*����x����GL6޲X&��ȪC�f��j6p�����FjD�ڜ'�t��S��JJ��O�`_i�kul���5\u&{u���Qo����1Rg�0mVO�� F�sO��6��WQ�jW�^c[(Y�6˱4!����̺�}���WkNM(�
^���<x� �q�$1`��@�;��d��8�.E��;[���t��7:��*��'��#vD+�XEE���u���o�ݲ]��H���'%x�:$�p�m�06��gYh�o����y�Ԫ��Ґ��(]�΄�.gܖ;������ׅ��zd����]�!�`hr2����}˒0X����cڠ>(����U������0������8����%%gr7'CT�� D�:�M`�n���B���W%>��SM�Z��"�[8����Ĭ�ri�ٴo�����^�a�}Խ�*лt�`ƕ���m.:S@��(>*�D!�/�\��ƻ��TB�oo\��^���/�*��Č�2��´_0�����#��&�rUm�r=�X�mOZ��.�a�G���:��Q��Z��獰����6��Q�d�鱩��:��&�Ǐ���WH�~�-�r�z��H�%�&g��5����Tݒ�����*��c����缐z܀Mn����r�@@xʗ�d��2<.r��9˱������mf�!�Ɂx��]��͈s�9�0�]1��"� d0aL�k
&���J��(�U�H `����K���g�� 0j��jmm��~9��t�]�~���a3~&0p�N���o#��P/��H|��4��O��tu�,G�X�����R�PC��i1��p��4"�3��$%�CC,��ׯ�]�s��������C���-�PC��Nn�#ڻ��%�Y��7�.�M��:A���sċ-�>}�/���T_�u���k"�C�<�g\o������ram��5��C�/����o�Ex�nkhh�|�:02�[:ܠ����uh1Wo�b��j�� ׬1bn� p�F �B)h.T�܉�xA�@@,aA?2�Nw�5�%���^�>N�`����8Ghh�j�� ��!�]`�(S�3S9���w�׏����fq�R"�)�:�_	##o?�ց��mYI�1��Lr���0ĬH����	+]��0���O�H�&�~���H��ӻ�}��y!�����@W�������ۿ�ۜk����ȑ����yyK�,�U�;�Z�2��/d�)�$#0���@�X��Je^lF�d���� ��z�.� p,-��D�����e����Y$�6 ހ��w'��A����ېSYY�05LE/����u�.��_�|�~�������0)�N2����RB�"���Xw1q�Sօ��=i��K�3O�JlQ�S��)��-셓���3Ņ2#�;�=@~�R�2��{�qVL}Οh�8��ɿlW���h\�5���["��=x���zl|�9%$56:��d�@�Y�	bl��� y�Z��1����>�[q�����~~���#U�+Z�K�:�:B���TI_���1��rRz� �d<,"�#��ҟ�8A���x� ��J��m�	�� ��k6�2V����D%6!�?p��8�����G4�-]1gC]q��0Pޠ���Kݵ�f-���0�a^2� ��5��v�H�
��Z�n���g�֎�)���/W�h�n#� A:�Q�7���p%wO��i�i��W�e�'��w	s������^#�������hL9`��W�>a�!%~n���_���N���'���k_�C� �P��[G{I������`OU���� ����0�W�*�v�Oy�m�.�.�����$�����A�փ���t�m��ʣ+Cx�%���H�M����Y;���Y{o��������?�����jJ-��U���M)�^��,�n����܄<��FH@��������|�Zr����?�����1�Cx\0l��[� ߸Tݯ�������U!����kxnz-�%V)'V5/�)k��;X�� �ѵ���~�Bj�h�5�F�D�'AE./[g��&�5��@ٍH���D��{N{��`�����"Z�Z�i���h>��	��ar��������f�Cg��Cɉ4�r6D�S.��������i�H�'�o��q�B�D���^����1=;��`,Zjb��(P1��Δ
��w���A�*�����)�i�}O!@mJj�uU�3�у ���O ]]�d�:ұ�~_��Q��Чť%!�#)o�hE�ħ���M�D*�M)����o�~�z��y�P7ˮ�a-�ccЕ����P:|u�B�/~'��|��ˉ.��a�6E�r��::��Smdr��N��ۻ$��?b\p���Kx�LY���H��}Eհ��gFq��9�t�H�È�U��>�C�90�P�&���ob�`�cE�����r������4S�����c�*���l������#�=�=���n]Ā�JO�<���h;b^K4��M��n���E�~�JK�;rr�[bd��Z�I*�:�@59s�iH04���#�_�?t
�����_E_9F��q^W�����ǫF=bcW�Фl��/(Z[/��Z?��Xf^��Dc�g�Z�l�ix��3��L97_^Y[R���٨h<�����SO=���C��[�~WG`��<����6K��tP%ǁ�ʻ�⦧���f)�:&�p�%�1'��� ���А@y�3( 4��1qj�~�\�6kP\�¼c�\���@^A���̃�B�x�I`XbI|Z1�ڴsaK�ƭ�#F�;�7� ���{�_�A�:zR�	�ql Sn��+[�%F��c)��,ĉ�"�I��ib�5�QHz@�^�����O����Ǹ�h��l�=�&�|#�#ZQm��a?�b���ǽ[���h����[f (t�2�P���`��Ʋ�:jH�6�-���?�T�/Xr�9:�51������ˤzڂ7-@���K�䮑,p���"ZP_1�5L~qt�v�~�`��A�ݘ�U0�bg��g��@��}(AQ6 �uz���x�ϩ�)�leK$��^.'��h������%��Ռ��1C	����X�	4����I�B�=�߯/tm�"���P6��wy�Y��բ�D��5H�JLLLZ�o���hUa���&�
��3���Đ�W�o�h�+�G����n��)-8���@��-��7T���y Y_h��w�{��~O�QdpB��S�+Y�آ^??���h6�p�D*]J ~�Do��CgѠM�8µ�����!�=��ߠ����f�x���e{�"$���צ�ѷ��S��r�_Lv"��%�+�7;�oh�m��t�xc�ֽo� ���� |�����@6�K*����hi��m<๧�?���^I�^�j�����v'Hfm���D����Nfff��(�/ο�@`-hN�_�N��F�(�&�/W��p^E1�pQVL>��DT�� R;O)�P�x��
A��'��BD D�O��g+�v��DFxu�"+�?EG���C�4~���BXa!�e*�C{�TU_���&^i,v}�8Bg�4"�U~�<�ژ�J}OKpWB�<&il�8�h8�ڮȚ��jNd�������U�~��1E�3a&$F�"᪭���19�"M�3��	3���+.��ц���옗v	�c3�*<��U�����{���#�jL��%�%�C6�����6��j��+D�2a�}T#-�]-dj1M����Y|�����!�zkfڄlҩ�����bNB����Iָ.��Z��ۮ��<����d�]�1�/��ȯn�C����6���kʋ��|�\RNlQ>�H��W���0�B$����8I�O�w=:�!C���S��#0�j����w<!vހ/��ob/zxgb6��<��L4=a0;�8��|뢙�7h�ǖv�þ~��sO,*_�l`�ZiMI>C�^V<Zb�HI	�{J���uR�o��� lJ��bTN��������C��YZB
/��'L��o��� (K�1Q����'|FE)�|38l8PHj|x�8$.Ņ1~�H�#��x_��o��7����n?�oS�����_�����4,ͼ�&'5mC��j��I�ג��8k��C
 �4�K�I�+*�Q@b�͑�<�%���0JlS6�/~#�g`׵ ($$Cm�]/������aC�,���\zt�(�>*5�
>��|P�H� }?�A4F�;,S��T�p��շ��r̵����U��ۉ��n��dg?���K��@F<i�'	cdt��q2 ���H8Q�K�lF��~���Z�A�a����[��<���lZ�՟*�;]�;���
���̩��+:��ɮ�)������h�/R�?���po<T6H��܎j+�Sb9D��p�z �r\� <$F.�C90��f��}�A*�G�Y��ܘx�H�V�8%o#u��~I��ΗeiQ$L>˳�L�<����")U�ٹol��D � >�~+�;���2�\ ��܄��7x.3�sF�@�6'����Ջ�'�een���Q�ɩ���Lo�*#���C��a�ÍZ��M�!��+����<��D�֣� Ji���|�x�]г����Ӵ����GF\ٮ��g�7Գ\/������Ѧ�<�ĕ,�T
�7
2�+���j���r�!?����A�a�Ļ��Ff��!]�y[$�_@Uv���󒏄W��dhi-^ B�Е�j�X�����p���˲�ϩV(g�{��r�������ld���p3�l�C��R3�h�&�5���u�L���K��Z�Y�w����k�$D���F:���1R��-W ��tFCC�]�7Q��: [�]��^�])?�߀<6>ؕ4[��R��:`D��� �w��}r��T�g�)�{9�6tB�M�9���b�!Կc��<G����@7��*<��\0��9��u�P�?v)�;p*`M|���+������4P��'�����O��6A�7A����<& ��l /�PSg���:͋q��T"f�dvZ�7�^<�f�B�}��N�h��-���&W@Bn���,?<G�T����f���N�i<ف7��%t�o�n)c��G�aVYW�P#:�j<	]Jy��F�Z=� �M��� ���ݨ1Q�`0�1�i��"\\*ܙIR���M�^�HJI$(B�f¨����"�)�S����E�O� ���8�բ
q��  ��t�ˊ��;b��G f����	���2
�O�`�X�s3тt�r2�.�֢G�ՏZ66@UVMU��%��\-�+���&,��![�b�vll��k�r��25���:{�芥�Bv�y��w ��M�y����^�]���4@}���#/��d vO�Ӑmྲྀ7����nnn���^?�g��d7 �����������7��s1�B}b��Ș���i6LB
j�C�� ��1�f��")�F�9T���1ZG�K�ٝ�b�t��������H}��cz��
{�d��f�{�%Ȇ���,�%����ᅊ>���.��� �ʹ,Ɵ�{��f!9O��]����pD\~1�#�q�hG�� ���>)1X�p� =�C�3����L].2�d�b����{�+�w ��m�"��/3��Q�������p���"�n�{�Q��w�s]�����DK/�Fb��B����)�b�p~�W�ϳ?��=.�����$r)�3p���q0ρ��H�O���.��lDmy���1}�)7B6D�R^�=7�G��s ƫH�&i�&x�0���Jv���y��[���E���2mT�F�i������gpY7���Y�C3=U�3��|3�%&:�v�ڪ'�7�STڑPi��ũ� �d~�-�=��[D/� �n�-���:��ބG!�\~��
���#��w���堁<ؗx�sa �-⓳�&q�X[ԭwI���@Ä���ld1�� !���dr4.�ԏiD[ ��)��g�Si_<=ۈ~��i�Zb�q�Ч��I���B<o��9�4d�Ү<%�M4Oi}���̞L1���ڑ�"���R�K�W�}\�yt����c���'Rw�t��<�Ҷ�M���zr��SSW��@Lj�8Y(֝����)���o�N�>��s��BH=˩-�o�L6$�+w߯�獴��٩�$j�~�!c��2��`���?��V�0�*"�'��� ��<s��U%�2��b�2
�AZ�Ԛ9�]2��eh+Y��f��)P�UZ������HHS��Vcv��8���� Oz�J�)��h�����-=ν�����nB.ń	����\�@=ٯQX����!��eL�iJp��;M�$$$�猛
���d� ��oȭ�^�h9>Wf�ۡl����L5�ݏG�)�25#�q�C�6��+��f#u��-�K?�(i��(���گǹ�Y?7O�q?���~�L�x��aw�	��dc�?@a0��C7VSs�F!�w1�����Zm%IH1k7���k��♏L[�؞\o{�Ԧ�Sџ��(�~���ȟ#:o���Xʭɛ�FO"��ҥK�?�0z��}\Q�����-�U!�����+?O����O�#f�9�Nȩ�"�pYcK�)p��c"��q�G	��tP8+++%w��p���s����@�X[[+5\��z9���*z��P6c�;-OPE���9�N�����d��H����>�����˝\Eu������ +��1�6�멹D7�O�@�BM߻�"�U��}����=g�/�ꛨII��gAg�s�h��ʼ��X�([ *��ny����f�U��Ǽ/�r+���2��_��2{n��!�=!��3�.��31{U�����sz�����'�����2\����$Mv���M��$��-�ꀿ��-�|F���D�)��V��X&��A��?�0K>B+0KrcH�=.����oX�B�ܟf���:�E�����1j��'�<uD:�^���P	�+��.����G�?񳶠R�A�րD
&�6�a�>]���Gd<iry��U2�ʻ��u}A}�fȵV��!׆so�@T|���n|]��)���lFkk�Q�����B��
E�ǫ��w�g������R=ryt�����ޱ� �I��ы�ܧ�C]�0�5n��:�f݊Y���mǾ��}ll4��- ��{9��ѓ��Ӗ�F�u�`���d��1 6d��
� �ۄӼ���g����e7��Rm74�F�.A��&p�U$�9����g-x�(�w&���N�E����`�TG{������x_��"���p0��]���G�r�D�ݵ�p�>y���A�om���s�N�[ԊX'\i�\?rTS�կv�2H@�X��.�f���k�����#�l�3������^
%	���E�����>�D��Sr�F��g��� ,����(��������O�"K�A�ӵ�V@�>Cں���?�-��Q�'!;��@���#��5:hM��	�}��g��,'Jd~��c�������_
tC&�.'�)���	�����e33JJ�G�㍏�_r��;��p�]c�?e{m3 JS �p����D���J� a��@�_3F֢��6v�6��������Ϝ >%桫�U�xKe�#G�V;ٯ�b�I<k�D7}qz��q��sj%���������X�+W�dH޻��Μ{� hɍ^��0�R�1[U�ͧ��q�P���'���b`��3>g͂�z�oɓx{�E}}�Ҁ�;}�[�.j9��}�km����w�f���&6�����V's�G]�xP��D���<\��o;U��]��!9����Lv��v����[e�+�o4���}�!�S�\��lE����g(�d
6%�?~,��+C)���'��-��󵩮��]Ko3�A���S��DT��Q������bѦ�"2�	wO��ē��a,���3a�#f�)J9���&�����A�f��΅�ׯ_�?'X"�bxB�K���y�Z�7PnK��5����+s1Y��X]���{)`�<^'0�qp/��_0r����=�(�V���ݟ�i��q=���7(I��c����pw-ޠ3�k�v����>~� s�d�BNT�K���4�{=#�3E���TWdP�)^�w��w[�C��K��X���I|�;�Aҭ@O�X~��vݿ��r���s�6bR�]�a��F���:�#&X�'����qG�RXҬ#Rr1��Q���(he�));i�5��q�kޖ�R���h����[A�]���� ~jqڸ���Z|5#�[?T�HO3w*�l�V��6By���3�)o:[BW�om俼ə�܄�	�U&�j%J��.�bTg��un���R2�=��۷oY���l:��[R�Eﮍ=�ä�u���96!�}��(��}q^����{�k�{ON��b,�&-wl���7���e����{���y��D*��x����M���V�լ�F�5H�Q(�����"�V�����T3�"[!)W�ZZ���K�G�D���@��~�B�n��T6��CRR���p�ѡ(����(|���/pa^��0e���mxEo4�H��j������Y���+g�ҼId������Q�����,��W���9S�,��-��g�3�T��J�)��*]}����!Apq�s����Ϳ�c���Z�|)�|i�(����&:�s�,��²�7J=��eW���ݎ����}��߱W�6�����A �&h�6����X�!*<l��.�'�S>���rc��܏�lB��IO�=����D����a<�z@������ӑ��&�H+@�ThӇ���[&�RD�8J}$YG�<Оy~������=��J��/��qy�q���J���6]}#�u1�|�$�T���	5�'&ބ�`<ˊ��Mx���ڜ�G�!�T	,�����O$���7�1hΐ�_��T��*=a9���+x�� �2vȈ~����Z�Rut�8��B���E������'��}lP�N懺S��G�؎pL�;�u�Ol|�����A��7���v	hh��(]��c`�	6$����9���%NjrU7���B^��7OU~��qN�'hOftƀ�̪>����]h�N�;�6���F<�e�rf��*���0ʌfh)�w�R\�¢RH�$�q.�Qʸ!-'�|z{(��3���6A���F��'��Oz���z)5���K � '�YJ-��;8\U$`�?��Ml����ZR�K�<}D MN�i(lxX�`S�y��`�`̀���Qu;�f�i<��Z�H������~7"<|r���]�3�E#�}TK�`��[��⁷pt��4�b��i�H��.q�����(Qڥ�0 ��r��1��C�����:Gf�'������S����R��O13e�/Hf�����+��/u�G�%8��xυ27f�@�tmrU�7{Xh!��0�,T������<��Vǅ�����Ȏ\(�zC���`e�y�O|���V�矶)ڲ3ߵ�k�Kwؾ`T�/�#��H��}�3����� �F�0x�>�:Ǚ�u}x�G-nM�Y�8G���c���|@�D#�In�/�zT/�*�R�DW��:'�_9�fڗ"d{?�n�S��tݟ�-=�R��������J����(T�aL�q<��r�� ��`*.�b��(F�-Ne�������Z�~������)���T���_&��i]�ϔ]��t� ���]�(
�����Ng�S��<f�Ԗˉ��o�̊�<�����T���rd������>���|��4ہ)l,�1T:��P2d�Lp�}8̧���'�)��Dm����`a�m�s=?N`;��V?��tCSE`=��K��2��Z�-\/�`�GZZX��U�{��%4���Mx75���G���eB��_���a�Ӎ"*ė�,�MR9�{�=�ɇ�_�f�����=��� ��p�?�s䨇}���׬�\��Q]Bm���A���J�W�c	�(��p��wa�Ú�8�-�L�bצC��W�\^�
ag�ߋ]���ͽ�D\�[��{���#���o�ǩC����7�8�tN��k*k/ m�d�H��dPs�*mH�B�H�6�χ�߯�uK�=��Xiz[��c-�6-���o�O���n�G�E����Pl���؅ �f���c��<|/��Ҥ�=��&;��͆����yl<j�뽵�������۵3���{B�03#���3��h�rhĵ=HA��f��)n�޻���b�uo2._���n>�_�5H�QW��C4v՚�8U�wQ/�9EΫA�_2Gsd��~l�_a V}%���8���#w����@t3�^��7�]%�5;�H^�b��3����'�y`~>s�l��FF���#�HǑ'F���p;��5c��o*�1Psˊ|� ͅ� �+c��'�@EtØ%�n��Y_�ڭ�Eaa�R!]��Y72�/ad��aέֺI��1��T�����o��^�i���x�%BY�s4��b�*�q�*$��A����jQ�|�;����'�0V~�!:��s�����)4Y��հ�6�Kgv5��_����c2N�WW�c���S7�d���}񹔆��\M��*�I�Zq�w8%�=&iߧ�?�&�w`��R�e���XA�|Sx������|�]c]o|��/�.��ϜP��ߢП�gԌ��~�m�=��߶�R��]���ӟ���"��x�:��|<����'iy�(48������]��������7��&����
�AbUX1��Y`�=���!�^3�v]�SB�?bD(�&a(�uf!���Vc�+j��a3�H5���U	P��l�p��7�'���|VXHڃc._ׄT��_;y��	��[�%�c-
�}Hۈ	�/HwN%d%�N���0�q�`�y��NK%�e��v����N���<{�����#2q�?�-Fsb@U��(�#�@����}���l����ۜ�n�O�	x*���%yfk�֬�Z���Ϩ�� �*78�Îb�<Z��i_Ȩ��h������k���8�Fq��3`��=Y���p�����R0��갚�ḃy
�ˌ�]W�UT��'!�F$�.��.�!D��U�9.��R�@ڗ����|��
�|����Ӽ��_�>��{_6�nk���j���	�����:A�1���N��_ nK��=����9y����F`;�^`��Ⴔ�B���L�o���՗�4�$�O�s@q�뒵���ꍂZ�%±�0���K) t��WY���R�F��'����������,�t�f�gL��}ڬ��6�6�Є�)��E��
��U�6�8WE�}���au�����y��fMě�l4����/ƙ���QZ??QD��, 
���]���{�L�q�����>?���4v9X�ɝ9������SK��+n�x�a
�d�嫯)�`�r��4�2����˶�ҙ�@R�J����:���������~Bk��(��<��洮����ɯq7�%�vR	�3K4E�c��N��؃�<�U�!�=��M�/���U>9��w���:�|_瑟Y�J�y��l��pw�x���ȓw�M��&�q�~�k�B�����Z�^�m�T�3K�*2H���Z��N�9��u�;a0YN���8���s�s��¢n��J�ez4>}�q��ٿ9*N�xP���*��s�{wAe�byܾt��w��r�bk;m�G����wZ����/���Ο��R�_8x�V��V�q��Z|�N�K���=U�����/�S�oWEF�'"�X������̞Lw��|*ӥ)u�/2+Fq�ǫ!��}�ǽ�z�]�c��AU˺qK����ɒ��3ݱ��нR�u�}�π�7/���]���d�mՁq�c��-��=k��J�٫�5h� ���Y��r$TM+헿ךlƨ��=:����=U�"�n��Pem�p�
1B~�x#��Ke29齙�'��~�H,�V�Ԉ�m�D�	��e�_���Q��5��)�%���;�0�� (��d+����줯�K4E�0��S)�Ǜ���Sw��h����PoI�v��2��#{oI�ԫ���*�;����mh,'�;�S�n�F���lM����՝�ӖC�pVpPj}/Ų���$|a��(}C/'B�؈��OH�jﺾJ������G=0�3��Q��$�zz�]��,nN���R��f�Og������DLC�a��A�ԓ��̡�aȡ��&]����C�� R�����}^��#�����Vg��~Tw��W__K�V�`'�?�>�*r�%���n�M<���p[$��w2?`�7E�zb��`�|�������5P�	��l���bu׷A9���/�$�?cʡ�u�^(~%m-o��6��������%Ѫ�8F$p��*$�|18)h�_�g�Jav��C�Vi~J.vR��7f*_�G�su��ڻ`����s��/��
�|1���*���Q���@�k�T؍��TW�p�W��g����?mP>�`z�y�Gڐ@B�_巣`4���Qۃ�Z�;�-:�1/z1��p�S����JPK%�$�!�������������>���M�W �F߸�����ӡYS���%���":7]�~���>�f찥��3D,����ٰ,p�,@s��`��_/�Vc��%����U��a���Bs��Էa�r�d�c��絭�#�F��L�ۧ��G�2F���
-� u�}a��<�P|g,|AH�!�Ɣij���6��ĉ��V$��]��<6�.7 *��N>��k[�c5,"�u�n`��<5�!5�o�����<d���z�R����P|��8�Ɲ�0���N��$��Q>��z�&.�o/߈�Rئ�'�d,�u�>H+���бƮ$�����^>cC�m̔k��p������U-�,x�L��b��q���o�A?g�������юh���,=3�'`��<��O�ϝ+E��J�,�+[{|�������V��xNF����Gm@����`u�X��o�)�m�����&�P_�,���`�9/C�=�g|ݸN^C�������*�-9.,9$��,������W��OE0Vc��n��k��4 �ԓ/��	&��X,�W�*�r���뻗8�oYG랉A��UBB��V-�#����˜��S_Ɠ��oS�)AH'���Ig�b���O�������`�l���;r�7Ի�:����m�m�:V�jQ@"�ٌ���j��UJ?>n<\Q�wy�X9�|�&��)4�!��2!mw����fO�G��}�����UC��Coķh��Q�mhj���[��s��)`��N�tӗż� �s��OFE�9p�:(�������l_{=�F�?{���_�<�s=s����j��&���R,�#��s��6�ثAM�FEk���"(��*p�p�1��~0�7+d\a���u���������p���*kڂ(5��m��J�3�#"~��?~o�k���ŹXP�Kŀ�Vc���V�fm@���'���Մ�u�@LK��R>�XԻ<*�$Zm��pX�5T��ߢ'm��y��w�B�1�k��²��⓲�ǯE$DN�f���7K
˸���{[/���6�ɝ�����om5��6tⵌ�Dm��*'�K�ޮ���jA�0�P�Ju7�,��;Nq����P�a7,��ȖA�Oٻ�啘�i�32.�����;z��E1U���]X	��������0~7u��N��2�*��{���A1�?o7d���z������v�/�;�h+���-DՌ�"�ޡ�\IG�Ϙ�)�O�j�U7<�j��@K�R!������T'�R�-�������X%�D��][�����ӭX�T4��Y�/�M误u䏓Q�>o^�U��X��vS��h��~���I�`Rt�w�g�͈���Y�����/#�3ƿ��wMx�1Z�����nCF�U�9p	k�=���Zc�Qܺ���ZtR��v�:}Cl��d��4��^_]�Ή����D��2��?s*���֭�Q��9{;l(R��Y�����#L~��P�\��1���%}���c��+�c;:	����/�vm�<d|vC�(O�8�t��˪�&���!���(��B���>�"���;$8흩X��Ŕh�缉޳�C�;�Y�g�p�D���G��V�������O�uy嘘�:,i�׼�䓊�bAz��6�ڿ;84����6�=�*��D>~�c��d&��p�.��P��a���r�U�!~�eͫOi���5Kb������CY0P+�[I��B������_=�U���*i��o�|�pV$���º�L�b5)�Z8Q�4�Vu�z�f�8]u�*�q\JP��J�*�}�0�\K�O0�~��P�����O �qY����o�W+��i_�ܜ���:{ ��mүуL�P�Tx�>�]�0�s�Uf�P9��;�����=��SS�|����r�Λ_�&����&�۞�]�]�l���,�z��C��ɒ��� �͐g��C[_����X��{�J���k��rwN�&�6ė	*��n��A"J�Z#��os7���jy���\�t�:�c��_d���U�-���Qo��fjLP����U�XA4+[�q�Y��b~�����qa��'2h�Ġ�ܻg�e���lY=EA�2����F-{�lZ��l���������w�_R�1�3��>%!�6SE�"��ƹ1���ua�>�xːü�_�3�-;��s%4w͑��1������P�n�}�CJ#~�1���R�E�;�>5Ξ�n}��q��"eK˄�eF�͛�Q~���bU�^���/�:ho�u�p|�w��zk�E���q�a'qO���ɬIcnQ?����"��q]3��R�)l�U�׈%�hD�����V��L�z5�ŧ� ����WC�pZN�gN�М�g���R��ɭ(Y��ΗP�_Z\%.�|"ehV�ST�t8׭��5���~��\��GI�����:�_���Lk'�-�LP>z\ɖ�9ob�D`��/ף2�T��9�:�h�=��ـp���e�z�n������h�T�G��T6�q�̞HY@���jo\���}�����Cv��d�x�.�d%1��S/OK54�$�����G��3�\����.x��y��ͽA�Y��w ��ֲ��US.�D��s�f�?���X�;=����o�0��	��׈&��F�����N�T����@�2�NRt����͡����/)��9s�
��&��Q�u�ǽ��(��l�8��t|��k7��������]��_���ؚɂ%�b/�z?�x���5�'9ƞ��w�N��6n֬;�FZ�Dd��\,�)���ʠeP�O�����^%��SCbڜZ�`m~���r\Q�(.��l`�b�91�8���P<$%q*fz����G���>��QB�*D^q,�M��<�$~���ɇ��R�D&��t_�ת l�2�����mQT)ۅ�u�K�e`AUtQ��б�χ�M���wR<}������u�tZ�[+��
��s�JJ��D"�r�?�0s��{�>^�/���|���,^��(�{y�?���F�H�M������I!���������\�i�h����*��;����N���(Rk�'��a��_��0ń�Ft��t|�8��gz�V)����(�aa^3��mt�L�����]��B��U?1�-���#��%�PoY}�{��6�cOQ�/�41�f�Ǧ�ecg��l�>2j�Z;i?��WqǓx���'ٵL<� �U�e+�1J�K�T���R�;D�Ƞ)-��wF�Z+U\,eMd֏4�_8MV�)o��o�m��� |��!2��ߒ)C;eP�®�k�[m,�T�)3�V�6�?>�y6�3vA���;���܅�ѥ��*�8�^�5V���{�;��K�	zП�n��u��y025���/V6HvƿQYu�����C弟�`N����1K������,I<9���|�z�����w�a�(1�ŭ���vy�d����]o�'R�`�k]X%V��%�JQgn	�#��U����N�l�����ܢ�ء�<�JfE����,��L��"�h�EW��@���9�pNe�.Z�j65�ٖ����:�I�R�����b�ȱ�����[���O�ڤ��y�L���E�~���,�h�N�N���PR�{��Ĉ�`������Y���7��qUV��{w
b~jr�
���u��-�i�:�9d�.)��+����eۈNt���Vqvtnw��V�3F�u�=m`N���Z#��|�7\�[��`�X>͇yWMl��0V�9l����t�M�g�r��ʨ��O���0'�)W�j��v��\��M���V�/�(��<ȃ$M�Мq�ʥr�%�U'�s@�%��ѣ݀�elˏn��,9.V7�z�S~L*��O�_ �N׌vo^+5Aw1�k���#yS���wh6���	�9_�ԕ\�u�$��o 7��I5���GQ����+ 9�QrO��ڟ	hH�}��/��\��x��2o�� ��i	��j?d�u���X��%!ɚ��c�p���>s���En�0��$8N�=�M��k�[��T��>�쥈��×
��m]�)~�H��ȑ�~�b1O��:˱�����>X��8����������lf ���{ϰ(� \E�EPTT�
"�!LdQ���$�!��dA@�"   9*I�HF���3[���{���{w/�9g`���ꪷު���\&�ڦ��������~��˹��
�'���W8�O�RE�ei�tI�ı��]��g��ʝ��^e�g)ݫr��+��gq�d��%@�C-����5���n:�|�+W�MC�BSV~hI��+6B��@���%���A��Ky�'�+||��~ϟ�^�ksJd�d{z�D%z{�'O����[�-y/L'Vx��2�P�-�y�}��,Ǵߵ���6�4H5Tb���L�$ne���b�Z$�{3R+I!�z�����'�m��UV������ Ý���u��S3�nʞܬGq��Z5�M܏U�5����%��W|�`�v��<n�����薈k���}_��W�3S��<P6����d�VVi� ���m��.��=����h,�����S��W�B�OP;�`lmCU����뫻W�i���lJM�5�уC�ɿ5�y��gR3|�����+�f�����3\[�?ݳ�=r�}���������']/)���[�fh���Ҩ�M���SO���[��h�W��� ���a%٥lǕKvo�V�P}|������k��n<2�U��S?W��s�����V����'Nd�o> ��(��[g��K�9�L_�2���-H$���S�e��i�J�9nm��F���<��%�W^��\���\z֢z��}�=�IA�{雗��!��
�6����Q�z(7��5Z2\�bR���M����w���X��	�Hާr>��+c�ƭ��L >t��FM�`�E��^�k���_G���J��zs�rd �7��-�Z�Oj�4[�<�yJ�����V�Xu�n��m��ʢ��ql�-"����FW����7�טZ�,�5�,�FƖ���g(��nm�z��=9*}C��<��'�i��mO���di�Bj�q,%т9o	��v��_}�"�JhD}`�_��t0�|S�"[��&� �>�+��W�S歼�C�s��2ç=���q��h�+;!�m�����r�����I6�����X��Ӣ�OE���|`����͂ڝ�RKL3$���O�
��Szn�ޓ!�ם"��[�[S~O��%H�ɋc��'�N
_�M��Y�t�|U~N�]�߉j��;3Gy�;�Rۑ�� [�K�7�6�A�%eu?���h	���^n�:'�5���#�3��+j�4x�F���GG ń��+�5�O8.���������k�o��D2�{�E|g���{wi���,4~����y ��� ��:��/χ L7\�7����J���3|K�D�5ǹ�Ж�gT|�z���x��hZy^�0�Ǚ�u�=��o��~�n@p�͎fhd�j�56�h}�r(���7��}�fRʂ�Ck��e~o�++,}o���vxqP;��U�����ǹgߙ�O,׷����������N�;V%:n����8�asنr׾0���ë�[vd8�����.vd��u�E�K���1y��RH��.�ĩ���*��7<si������wr�I0��ZQ�ڼ���Ϲq���� ��[�4:�}N�[/z/��s�Ӊ�It�dN�*�n/�̻0�f�{O�]ɍ�����
��D��-[6f�F��2��?�>V��'��NX��$�(s�ߥLz�=l�<�6f��#~׾/����zG<|4b�\=�E
]��Ќ���<|�b����Sz������a�ƽ��_9�}����bQ�ѦS7�͟�S�h�;e7I��v��;�O���^J����o�K���͙'�]X��+���?���S.�����H�:�w%��;4J8Q�?y�|���ע�!�&X�Lh�o[!?P�lq�C�Oݏӹ�'�D�}J�9=��</}e���w���}O�};rY�e]�3��l0��Q����}�ޘךϔ�KZkr���Nq2�_z�p,�߲���,�������	'�H��>�]s}��9��[����W��W��On��sU�n&m�������:�g�K.�,VtF{�*01�-Ŝ^C�Z�ރ��5�oH���O�V��t�|�ؒ�woU�>�c��?]J&�=��d��|q�pCV��v������_�z�L�U����l7��&�]�!%ٝ~_�������+�ϾԴ[5�mE5`���뗛��ľo?�m��Ή�į�*?����۱:xF�髯��"����Jc�e���ON�#�������}ږMۙ<n�\:yl#��MΒ�y�?]�,f�1��ʱ͗_��sYS��_1��s�(�۶���fP�N~�4L5��V]�RH,�7,<�����F�&���I��w���AJ�geVӺ:�퇍i½F
�%
Dw$�7��(��c�"M�;�%
��sVT�Z,pqCyKsó�;�N�J�Q�
��J&1�<m�*QN����#�t�~Z������[ڛl��Ժ�R��9���3�c�����LVsg���5�=V���:h|"��zL<I�?X7H�~JpLs�̴\hg>4d�h��3Y����K	��{(a�E���M�6�#��b��	�ܶ��_�����J��H�*�����[2�.�ʝZ�d\�M��,�pƑr,����ˮ�+#�������{��������]|���A@E�5�F�hOE�81qo�b,�.>�k4�G9f��{�ݗC�
��R�:��D��S�i�GJ�56m9�1E�x�tT������7SRJ�x9��hIF����S'f����9T����b|�j�S������ܙ�./�/���O�s?8á��c�N��n͍r?����~����S"@a��]���ゃ��*�^`6���
�S�5\���F�sg�<�l�ݶ�j��
5)s�ۖ�z>��d��n�8��c��@���޸����.�d�"��9�C9��?��fi����J�Y8�{�&�J����9	�iŜ���#�&�<-�8���^����,��Plq�>�lyZ�~�H��Z�-�cm�6+�3�q�z1er��Q�Q�������D���T��kdJ�vf�>X��<�T/T)6\ju	��d*&���L9�;�30��ޮf�MC���mU]Z�!�J��}�-������Z��à�Z'�A�e��n�!1N�)�������� /L�9{�!!�^��3l�Y���.'ǩji��2�ތ��v����X�<�9�:��n����Ie7)�����Ws6H(�f����MY�Vs�¸���a�3�}�G���˴^�t�՚�/w����۟�2�,�qϲޜ�&�����|E��vYtC�n˔�)A��M-�-�5����H���]��`�i)~Gmqt7���;��2y��Ȼ�ߕe�Q�dO�u�p�гTt7����	�B�吗�����К������6*4&
W0u̴j��|籤��(I*u���>Q���+vw�^�u�mlc6�� �M�F)�������em݆��w�#��i�M�F��H��U����e�����FB~	^�����NL���j-�`Z����c���c&���6$��3L�LԪ���h/;LFv��z�}9}���g����$z7�*�פ���
�+��O������7�?�4r@�5e��m��N˦a2���]�?M���1�'�u@J���8Q#x�;[�}~�5�V뇅���WW��R����$u�:yTװ°yOot��^��-hL�<�n��M�Gh*��d��-n�[�Qy�o����>
�b0�ْ+4�B���@q.p�e�g�=����[�lI:����c��;9�i�bI�N;�l���������P�tQ4҃i��$oF��_'��~�uS�}���`&���Mf(��{;���P���gϲ߾��}�t��g�6?\X�L%=%Vkx�e��Ȝb2��r$W�s�G?H�ّ�2��W��'M��i`y����!�o?��3"��?������$��Ӣ"�5�R��]Ф��]-�nl�J=�k��̍�M��d3�:[�4�<�����Б$�7_���������<cf��V܆��P��3���C7Zw5��j�(`�f�d#�N�0{�Շ��֎�*��\��%�J�zu�GD�TFp2�Ns�VG\ԃ��־�c,e�������^�`������6�Qy��u	�_��Qޫ ����{��y�"y��*S�p	Ec��g����7������(�?!�yg�-�����ݯ�����+ct3[H-�Nw�>����^Pʗ��H\"MńgK3zn#<g��$�#��ډ�훇�=��2�6�����!\o��f����*+�����;]/^p�1L���53:���4Ϛ�:MZX�$�D�����	�C5�	�Ő�6�)I�_�A�~��&�~������;Z������I�؃j,#�:D����saN�V:9����ī��J��_�d�|Wj�2�>��mԈ�E]�~5�g��J�ͭ� E���j�ڷ��Bݐ�V�@�|�u�P�nv�k4�:H�)U��G�)�vɐ}��L�M��k�!)8�����st�;Ty����=)�3� �Q/�'V��^���gk��q�B�L����P������|�iG6l��oQZ&�~a����{����w��3Z��;��fw*�i�Kp�Շ�˯��ߋEI_����M��F-�]�v�)�mF*�Z���.�0�T����g��E;�?j���|cMgǴ�ˡ_�5��>E������o��Ye�33�H??���l�i��5�xp �)����?_�F��g*�g��rMp�;�Ln�d�2�MQ��z�&��|��Z8��ģ��ޟ���	;�w����ۆ|`�ܞ�J�d����E�]�_��N��o�������]^�.�O��'h�z��X��u��"�E��\�.r]��U�+Uq���|�xjP�g��G�{~�����O��?�Z���i�����O��?�Z���i�����_rjLL���Y8�q�s{���[g�Pܣ,xGⱑ��wS��iՅ�މ��ֺqqI&{k*=��:��w��S��������T����x�ߒ��~����,��������u����\�.p]��u������U�G�	�#�b��ȓ>~��ӄ�F���1S6	�o�"�����y�>��t?��(&�md��]����2�8,���L4,Mx��Г�ݽ83S��}Bȫ��S�P�|7�͓��V�D�i�H�Ȭ�Z�xTEO��e��,6MU6J����2U�`J��l��ϯ�eU�.p]��,0�?��]6��5��3��RV�%�Wv�;,�\�������̛%�/�g�_�5�1]֤>�g��1�ǉy�B�sU��|��ݨ��v�8���#}�������Y�����br����ݪ|�̌q��k\�.r]��u��"�E��\�.r]��u��"������ �o��gb���Lmm����Jm]�%{������a[��Xm}}����B�b��*�鮮����\	�� .��� .JJ���>~�~�7B�g���.Z�k^����7 i�E�8w�N�g��[{<<<�~~�/�����+./_3�0??��cPa���Ϙ�(� TTT���虐�p��A75����t0��9�����c�߬�����ի��������ׯ���	��(��������S��TWW��:p��0Hx1x0Ix|~��k�g��h��ٟ�;��6 ����64�c�>��~JN�dkk�)�>~M}�%�RU�16߫�||fff�x|���,�4)O/hβ�A�@����`{��A�F�mҮ`�dɻ���X��U����xCMMm�×l��zz.h13m�LG;[��LgG6fZ����[�.�|����Naئ.�677���:WVV����4J;r��\uһ�����V77�y	�_s��(l˶�
4�qiʹ,N�(ަJz������6G+�%�oJDC��i�_�	���6h�52���mc�\�|�zC�J���0�Iǹ78˸^�ձ�E�8�=�N�Ŵ�P�z�ko_�K�Y�~a=q߫����9Ϝ�S���f$l�^$��*���F2���;������LNM]266V6-�wI��XwE ���Ru{;�NU���쯗ҝ1�9��˳�֤�������bѠ��jN��ąߎ�/�"*{3<3���ٕ���Ƒ3{Tda0�1�XVJ-LzI��A��(4K�o%iK~������c��Yk�E�Qk2Zi�%n�p����%i��;���'t�PʹZ�M��W�+Oҳ{�f�:]�;Ǌ�T2�[���������E�|we7ڣ3]����08����}�+�|�����HfOz��8�aw/�ypL�I���;���8�v��0r�`�綱�Wf�~v�|(������ܯ�cs=���C?��O��_}xT{X/V.J,Vh�Q���Mu�~�Myy*��8p�?5�;�F#�+9�����9b0V#����{R���J��A�R����;ev	d�SS����`w�s�����
ܙ�ƽ�lmm����000�6��Ps�I�#��->w9��ʪ�3���B�.IKKM��'��}�9���Z���M���y(�Z�uHPa�����M��1�XĦ}�&�)5�F��^�����lPs�<����N�3u���D�#�@�g�/^����l�cӕ���_/���r���$�R�ӥ��m��$iW�N4���S�u�x��2�\!

���ݢ�q$u�)_��:|����:Щ��S��[�8Um��hU��
�ۼ{�K��D�U�@��/O����XJ-��9x������0�Ϋ���p�̞is�M�/�Y}z�����@~~�i�$�>aR�y�����:E�C�<�B+����-a=y�5�>� >���f̥*x�aa/B�ͷ���vGQ�F� r�h����;�[Y�e�������9@R��?������W�up�r��������E���B�-����Ѐ��{��"�6�܌A��3��%�%��m�l��K�Sc݁�E<����09M�c�8�T'I��{�޹P����~j�����n�t��]O�I)��;�S��F�!ŹRX5���l��v�v{�j���6��h> ����۪h��w���?^WSCe�=u��0��mߩ�.��.Dʫy')+/3������a�f�,((�D��(L/W�cojty�]����׵�/f���$�L��E�~��m׽`Gr��gQ�܌e�ٶ薍ۙ�xf"�>�bͅ2��M�g�n*�,��aQ�U�/�� ��5ި�}/��\/��լ)�<��}%ZN�%JS���{�^-YY��'{����yfݞU"FE=�^%Peq�����~lz}f�UKz��U�I�<bo�J*I֔���i2�S���/w�ªu@Տ���^�����ʤ4���["(��d���0ĩ_�~���ɉ�*�;��<����[�@���U��l7;
_��C��i7d��v�1�֚�TΠM�)T�!�S[�o����H�L�n��lsC����vUH�fnN�Ѓ�O��M�T�����Ӹ�t_��J�����/؛��h��S��~�	KN��ne~��}�>U}�1��u��ϋ�/���ܯ�<�����:��-���E�~��=�2zʗ�Ҟ@���:��J&q͵��܁L%��k������A���wg��g�s��ͮ�Io��.�ğ�*��2�4����e#s���}r����eذ����.�P����GJ�7��I�
�lŷ�$��N�|H�d��@��[�K�DO
���:��{�awF��fy�WY�#2��^�mMK�b�>=h䬔���s.J���fө:E���Ϣ�T}1�3�m���O[��
��i�%�?��D����A)��1��]<��ͷr.������k
�݇��-���ݰY��~]<��(�L����8����Л�n=�[2 �w��st��9JcnaQ1�q��݁)� 0S	SR&X��!6&&�H�k�>}�$����tT�[�y������8�{�bǁ��+��x�F;f��r�U,nd�~��D�N����%D�_�CM�rvn̰0@�l�˫�JZ��Jh����� ��>UZ\jJJѷЋ��e9�Z���g�W�e��/]sS;��h�X!���������xR�COy�PP��|C�H��t�����奅�.���0؍~nL3�+�B����Tc������T ������_s���|M-���2u��v�3�ť�{����_׼�	s-+%v�/��+Y<h��8�c���pQ[�WL0�*�R<_{���tg½���+���v{qU�3U�F��gZ�4`B.O*F��8� S��������������0����{m��������� �3#UR���B��Ϯ| R��A� LT��J	�Ef���^�S�7i!R��2�a֨�▆{�5�ű[i&������3t+o�A%�7gy*��������N#>x��T����S ��Jݠl&ini�g�m�.Q�E�mA���75�:tȴ�`Y�'��;""�F-V�GV�ԁS�kW�������$��eO7ϖ*�xH!)�5�NO	��Τ���(A���3��n4�K3:=��[v@�ޔ���˪}���v5�bl�
�H`�≛q��v-Do���]�[��Ew�!�
r�����ٹ*G��ed]������N���u��ҿ�{�8�HU!$4~����X����%����o������
^�n2����:ؒΕ3�a\PH�F�,+x%.��N!~���*q�hk��X�,���9�KDx�xx�bX�g{�)���O����R@zh7b��v�#�Bc0"�x�|H`��m��I)m�:�A�e��:,��?M���N�x�������w�oލ�9����Y�,�3�M$��Un}x�G_��hG���EE��*-�u�}hT������b@�^J������q.��/Q�8��)���W{�oOň�瑟�A��񘋴X��}�<]Qg�[ס+	l���=>��ZG,���5#��k�E���<-5I��w�\��;s��M�ԇ��vghR⒳��Ei!5*�d}K�YE�.��*v6�WT����wZ�8M��vק��������J�����d����-�=q���~)k�~�m�ɛ���� X�|mꢽV!{��JA�7s�� c����e��vl= ɢ9~��]�N���(m�;�l��2�@>R�#5{Ȱ�vu�QZ@�sWv�%c�|��𸡶lfٖ9��u�MY�Bf+:_���z2ι���.2NŬ��Ӽ�� �M��I(
�D��.Ͽ��tu��Mo�l`�\�d��m�:�%=N�g�}u��+�\*�.�HIkf��Tٌ��7���yN�bQV����1���-������b�W��TLuM�K��_��;�+/�V����VU���J9I\���`fG��ҫ��4�fm��0<R�h��0�N\�BL�lc�H��(T{�]�i[񯒗0�w����|����"M�h��-�&ʹ�X-t:\�J$m��7��!t*C&;�w�}Vܮ�^R��O38��P���D5�'c �A��#������h-�ތ)�]��[xȲ��Gc�����%��<rC"�������ۗc�o��pRU��$�~yJm�'geiD'�~��P���!�6qo�򸼔���egl!�F� ��WIJ���Lt��b3�*����0��r|�u��`f ��`�9 *��w��)��4�R�� '�;
;��Y�"ӻ��R�"WE��g�۲��"`���T,[����K�<���Q��^��y���N���P�R@����=��J;��`�s��~a����{��Q�f��kF�����6\:��[�Nh��>9�����s��JP%��������^�u��寉!22�t���B�Q�M<	U-@<�
���|�e�㭳c]]����$y;&^���ug��� �q���s�A^M��V:ƹ��t������kz�y�v�;�9�^�u~��{,8����B���޾��+<���4@�$��`��.>��� ��Dۇ�� ��J5�~�WV^���*:?����]�\0�{i3؎*�M�Q�ɞ���f�7���X���o�%q�y0vW�SE�NI�>�cjEح\{<��00~�#�E�4�W��N!'[���Z�N$uQe������
�Ri7��^Q���/*�N@�8����Rǵ+��I�B��1��Z����dM�����J��������:��eI��d���,���{R��T��a�1*�%r��3��8z���/h��g���l�%�m��ݹQ��q�0�1�bL]�@#W�L�Vd�i�j��i����P&j��	��({���B!�Xz�=�~�m�U� .�"H��P������`,,1U4'h�}�D���v$�02XS'R��a�\����91'Ǘ͊;"{K��f�H�@u��2wA/�;��z�6	�d���혧`�{]c���I&?��J5ė�E��I>��.���r����΍ahq����Cy�E'̱�xGP̉����>i����!cG[��Uq!rB!0��*戹�*���Ҳʐ�V��رr�*Mj#�I���W1��:�iy�`Rl�UK�by��֐I��fMF�I�r���7�m�թ���Ԣ@�:Ss����:��%��?Q��jɣC6�,�b��)�b��<d6Q�WiA׶�W��[��"c���Rx�Ĺ�?�{R欗��-;�WU�,-���W����@{��t"f�V�7]��Ѿn����2依=��ږ�� w��pKz�VV�M n~�������>V�6[ħͼ*��/lYo�ԡ30�Ŏ-M[}Z�!�'rm���)z/�f�������TȀ ;t͏<����`7,
��e�ܹmܜ�1߭�����<�2x�|;���~U���V,�j�P�����3�$ˤX�c��!4ю�jev��*�����4.��� :u}��*���;.̂�6䦂��/ʞ�6H���>�|皟
$Ȧ/�bn�:ʜ��:��L��2��k�Ɛ`�~�'���O �*{���|+�����h~�Z~���A¸��!�^x�N�}�, pX3�?1�>ɀ|�t/`�vz��s����W���	d��@�"ޡ�]�UYH���[OHR��I��⡂8��THJ���!R �{�.PE����hs�%�t�K�X�y��!�VP�ؗ� U.q��Vu۩�=�
ZP��)~��%�kc5��ܸ�3\��X��G����s8�}�w���Pk&_�%�E�~I���NNN�T���Sa�FaV�)��>�Kj�@���:����H����8A�8��_%0�������˶ ���R���\��?��S����}2igU��	��?��K�uvX�/�y�'j�Ĩ�|��H�;K���+��҈�A�����&���VL��Q|��ҡ���]��o�b�,D:�j���`�T�?���W��rQ����d����mY�_�ì6�S���)���0�0SW��뫫_�ri��5�|�i};r�z*QIO�������v�+֬J���Pq�|U6pv����[�+Y
�0�����P�g"~�#�v�0Þ�fX4m5iO1�`^��[���n�Xd�)�x=#����L���_/��*@`��ǻa�Ϊ���ޞ�a^�:
�f�3��[$l����\�Ji^��,]���dMt��{�˫J��g`��%:�����:��8�@�gF]7"��c��xh�n"W��� ��}�G��^ù+˫��"�Y��p	�J��9�^ ��y������}��$o�
A�3�QYe��A𓸴NW��_u�d�`'_�s����� �
=��ӟ@\������9J�/�*�D�sdϴ�9�P1=?r1�k�rAA�D��׃E����ag(r�#����!�Xܥ�Оc�ը��_�iE�9�ҢJxF��:�vlQ_dp��l�C[�T,)$���F�,����[	GsH>�/�T�R2��%���a�79��A���.&�d\��ᩞ��=O�I��:qC�_!2�F��(�I2�qV�q��zZ������ TW)�e3-G<1+�V�d�ikֿ�n4:�fړ#�8���0Hp2��O����P��6��|.�}�ɜ�zs ��+�#+�#��rK�P(#�c5���%Q}G��F��Rs1���3�h�JZ��,;��̫W����Yє�M{�D�u��ϪE>��\�3]+�щP��+�'Nlt˟q䥅}a�Μ�a7T�]�GJUHuG�X ��Mz�Z�&Z��E��`��m�#���섩�I�K�*�Q􍓮K3��S��o��*�ܤ����I�Q�$X8��uG�y�w,���ϴPi���rR5[Y�Ꜭ���x�TwTd���A> �|ƪ���Ӯ�B�w���?b�d�;P��;Z��
˃�zy�*�X
��]�����`V	���,��皶�9.�a<nu^���}� �� 6Ѝj�qqq�;zy�vxAz"�e<�N#{���2
�H�����Ӱ��P	j�+�<CګM���T(`p	����n_ �a)��|"��VT�ƒ?�\��x��B����� ��Taʫ<dV�	q�f�/2�*�!V%�e��d}�Y/��� *��ɒJ��3�ˋ0#~й}��o5��]à_P�3Bx��1��j�]��=K+;�����X@"��!�J�	���k9��,t��`F�g���W��SIh��m �92�"���������Ǖ%��R��'+U	��m[`}H�*p[Ѣ�*�S�����T�JƄ�A�GT���G�"��^��}��M��]}�y`���@=�Ѕ#��G��"5�ei@�a�A���d�o�BbP�Y����,�	\C�HW�����'�AQgM"O�.�`N���(��\��D �+]~.�~w�_0ѯ|��d�`{��X
����aT�����Ɯ��
f��zG.�)5�oZgzW�3R�Yv����4-�#m����b@��\Ǖ|F�x
���v�=�l�?�H�NÈ>s;):$S��e�D��j�fO��\�D���@m��Y\GG�j6��JBL'AgMەW��emT��*�����t0 �i�����Ge�y/`֍�m��Pe+'�^Ǫa�{h�G��	!`[_6���%Z��@��N/�������-��kpGR��lU��`�n�lx�Z���/��W��*԰d;�μ��3(E"f�a������"Ff,>�E�a�o[�QصZ�.`���gF�	���qz����S��D>�#Яt�ݯ0=���U���j��o�M4Lg��@��☌�շ{5�=+*;�P�����9��o��K@i�Dl�rxNl����~uq~`��ZRM>Zc�L��9�ꅮ�0_�+��ܬ^�N������"��^C+��"��BEn�% �`�n���4X���YM\-!9]T�KF��?Q�D�j�.~#u��A# 䁴�\TrP�����RI�����`��2A.Dd�ΘCyN!*#,,�KKT6�3�w\���]�- gi��5"ՐW�Rk��o%j^!��6���������m�6�>�b�+���3Wj�l�@�۱�뭵?��^?� ,B��h���Q��tb~q3*��ٲ�
\�4&{��h���X)�H�t�JT�-u�h�$�����vt|~���ݹ�AWH91a�>n$��~�@\�����o��X�m"
��DſI+��}��;�aO��^x�`��U@?�I��ۧԚl��W���/7&h�Q��Lvzq�S�{�pZ�l�j9�]�)��zdSwQ��B(�	7R����":����W�*�	/��
��APS=�`)�P�Yl4]�cA�%�T��"���yZ���f���l�\j7�V��'�l��A���>���BZZ�A�0��K��w0SwC*P;��Lf;8��dMO�5DuzJXWx��~2��%1l ��~���=�b�(b��E�N���^�������PӏN�P�]�Θ]&�������#�k׮�r⮓π��c�$.~1���K�.�w�4p�#��O�f�l�Y��$�Q,��ɨ3�f��$�J?	��Ѩed��c8�]�k{{{���v=&�k�Ζ��?����>�p�T��J�/���;׃J��o{��� �Bd��լ�q�v1�Cd���Iim�J�6[�eY�<�Q<��-�b�N�}��s���аi����*&ƧP}����B2L�CI���ݺ�{��D�9! ��τD�����3E��	��fT�k�u����}WX���3RX6�'�H�~2�#������s�:���  KK����]��$.B�&�t`	��?l�8*PP�!D	=C1�S��t��D7���Vn�;)׽��"ĽeZ�<����>�����顐��^>��}��t�&� .mx���p���a�Lm�,iG6�F6j����;*����SJ�����' ���	��tU��o�b��˨'�/�m���k�>z���ն�U�]��Q���+!��f�C,ot<��{螘�G� ^� R;��@�n�yq
�
O�{�8}-��!����1C������fj��U�Ċ+q��-�����C�V�$`|�THxV���G_��h����V:�N)�ݲ��|��x>`�%��љ^�L�ӝ@/�<$ȍ5�҃`� QvȬ���5p�����y �9�VW�K\g��u��8]Xe��j^�o��S��@ǆ͟w�&�ο{����gZ�V34��Ds�6� z�;wrK����P_-��Rq>���p�b�२���R:��XQ�J���m�RQ������F����`Gb]B�����T>S{�Q��h��ÏpZ\0����R����L��O7��x��?}8�#�8�b�����N���C8�����D���c
��j܁���?u"���kѥ��.%<U:�/m$��y������o��?�M��<�ǠP���B��Tx2��蚘#���_d�RY�A=�� ��L���g�3L���}���T(_�t����~�5�����܈UJȈ�N��㶼rt���pSfXt�c��r5F�s��7~��~ ���j�4��Lf?V�##2���E���P�Ox渲ܴ��p��[���Rr?O�E@��S��Vߐ�sC[?BE|f��͖�a�^���_eA��Q��O5�o-]�z@�+IaB�X���.��n��Lo������(E��8��(ۍ��h�'��t�^LQ�e��'N��)q2b��C�ܟ�K���X�;+��디��M���>(�4�+��j�UtDP��6v$Q�l^���b�s�zo`���u��n�tJT�e �p����c��� �Fg���͍X@[�Ȇx�=<�y�l�3��.�^�b�9u2��K3���%��,���yc���ym�%NH|�(�+�ؙOB�,���x��:V6w��:��dc�LW��Hd�c���
Ԕ)�ho�G�IЭ���1�U��##�e�8�|������2lQ籨*�jX�ܦ�X�M��B�� <����{�N�9�Wو!�c�o����AF$�!~9��1�1!���vz3.e�4o���N�6���EPU�3x#�#�����cJ�	�rD�����S��E�$_���d�>���߉�3��k7�(��uэ��D��b�9�4?�*�:���d���! U���'��b̏����`���
�%d,--O�I9�5^�F���v�ޓH( ���o�>T�n�����TYZ����h;�32o�����aM�j���{�S���,�&��3{�p�%��� �l�����O͙�m�j���=�c�t����5�a=�,�Ļ27s$)@߉(����E��ag0.�@�������بc糬;ZX���mo�W%li�D.��s��[�C�Cݱ/�$�;ܳm�l�U����q`J����W��������UR�HC�Q����/�e+�}q<� �W��m�Q~N�U��X����P�9"*;^�Z�c���#��OU��6�ӨC*ܶ�N���¼l�f�2����6�; P��A�PC��`77�����%�@�L�IÖ��@ �z�ԡ�.�xk�M�c�Jm�K}X����CҀ�a�>���7~	��b%�q[��&�m����bv�F��;��vgq�&u�<��+�0�L�J� 9��e��i��o�C䨙�an�I��ڹX�.��:���E��N��,��6:A��'�k	96�9b�:>�ժ��g�8M;wX]B݄8����*gM����3��t|8_axLuR1��JbC~H<�Î[��S�&�=������7�I.��~E�M�O�Kҩ��qQ��C�m�Qi��_���]ѡ�i���#�`l���|�.����V�P"�3�̛�z��^7d� ���$ v�f�m�~�\W�~�e�3��]!�հ�]K#@U�U�>g��N͏�� �o��v�p$"m .��q#�76G���A�g6(_�l_�4�.X�֕��Nv]�JBuC���?�N0�^}+���V��9�ٗ��g�u1��oXO0A��W�s�?U0���(B�u(*%5U���&ԡOܢ����f���:�Z�A��u�C�(2��K��x+,�5�&�>�Z;�|L�X?0��_���U�v!F�X�\H���8.�qj��-�B�B9.�HZ��.tq��S�ڂv�k_���'�?;G[vĬ8d=��ܹ
c ���$w/��O�zN�>�l���y�LP��+BJV��ٶ���Hݎ���d洚��#��6�x��6�m���^����3��!v2��P��EW;�D侳�x[�x���9��)�j/=��h����'4�a4qy�-|��nk��ßSCO�3��1�8#q(Q���{��0�`��D�B�Q�^R�b'u�|md"�*�n��6���A1M@�O |�#AC�Ųݞ䫇�4U��{�_�ӧO��Z4h�Ȩ�ԉ���џ�I�t�ۇ'Z�uʉԞ!�b@���Η�������h$���O+%F�j��M��F�'q�D�F��򀗄��;Z��~���ܬ�: h��w��Ϳ#i:��F��5�F�+�u�j�,��ǌ�q�^<��	Gp��b����:Z�>j��C�S$#���q��>~�Y{���~����-�=��;w`y7څdo^{u����`fF�o��tbJ�Ψs�V?��R��R�Fi����yԞ�A!�)��%���E෡��"k����iw $���
�pd ����w{*	��+�<<w��^Β�Ld2�_�L��e���y�L�v�/�Y]��	˖�R ���hy+�m�J*�3ˎ�N��o��5콳�E��m\��:����K�7
�>V�6("�d� �J_�U)o^�f}��ia�.'�~��(�;w��91Y��ڧ팑c��6��T�-,���~ZV�|�h�9�F��S���D��*u7L�~���o�NI-�iP~I��B���G`�Xs�2���_w�x[CK���X*
?"A�#L��r��%S+�.@���@����+��M�<@aޠ���"�w�(v3�Өٙ�)��}�[.��$޳�3�
�tՀ��s%҉\�QK��T�4���U��d��TJE������X����Xq���:OA�q�A>#��a}'�����n�rN돎�5�7�S�t��K�`�����9yO�ׄsވ�`�)ٴt�q�lQ׮:��b��O4�m
9�������l�U�Aw�р*��t �����N���7`�Z����,�
NyO��u<���`f�۵��~��'d#�ws�w;<'�P�
��8�o����-�d�8��K������޽��������� .�/�ϘtTΆ1�Z���5Ң�,e����젎h ��>������(�p����F���zh��~t�i �"����������p�xU�����ml>DA`2�D0A��C��m�;���0ӯ��^كZ��W%��R����Z��OqOzZ�׿V�|�J\���Z���<�m�#�vK�?�N:8揎0kD�^�A*��!�%Q�?LN���{�1pN��.&� ��Y��j��,[L���B|��+S��Αu�d~y��1r,���z -	xdc��4L���H8�]�Ī(�&���k�m&�E�!K1���ذv�O���|?R�a\�x�l}jξ�;K�Xw�[�{�3툧�D�.?L5���������}���"����c*~j��r|C��E)9v����M�
����q��MmQ���[����!����ne-�������-��SAqea��站��<��ۙы�����P���4d\���_�ol<�y1Z�������b"�%]=�
وnƿ�K����x�Nf�u�~$�,3:���e�9�X:҄�{�J)��yC�z8�ͺ�K�XO�[=�^�������/2�;�:�D�1g��!Y��a�8<�j˿ՔM��Kxy��1m֋Ԋ����-���N%�'��S/�)������@�w�nǹA����sU��6L��6��~ԃ��m�/x��ۣ���@m�N��S���/U�����la,�'F1~5���nA�X����.Q�������{� �KA�U�sd��;�܅��@���xDM�q$�7o�*1��yᾛ�O��`bo��d�`s�I�ܥi�o���[��k{��]F7��,�g+&��?R�+���� ������� �A�X�a�7)&Ǯ,N���a5k�$<�6wu�q�3�3�����Vvz-�z��;�t�>���n�c�0ٴ��c'ԛ?�a�,��(�����G�tT�z�AB�ɸ���%L�'��R���%S���C�%�ǜ1�i�(���������6�����c��p����]@=>�Ÿ冲cE�T�Ie�7t�?(��0LEy���[#j��zN+k�K���[q'�MC(����?��������]�Y��Qx���S�j����<��p�梕9�f�� B� ���K���4.C� ؾ�	�2��{c&T^�{�kyaR(��'$]GW�)�)%Ȋ�C�d�`bY���c�$��}`�R,-��������Zv!?��^D/� ��-�r�ڣ���-��"���q���X|%j�.!H͂lzt��/je�o��400�����:$'GdU]ǯ�B��XS�:Z������"t�h�=��aqv��2�*x���3�Ti%�[��]
�z��UWn^^mfS�-֧��G;,WTT4m��;���S��sP����}D���
|���K�{_�s����X����2m��D��5�]B�)IѦU+c���l�B�U���	-%�G{J��}_�uݟ���u�;��:���<��x>�z��u�o�(v;쫌NH�s����A%0�x���)����t>Rń%0�B����	��������o�uvLo�����v@�����!b�]-�,9�6;����`��d�Js�n��k�u5%�e�3}W=fg��Jص�w*u���N�9�9�軿�x�@��� �k�,絳i�%VV�Y���=Qe#��0ծ�X���J�^�BG�|��ϯ�0�(ɛ]��>=1f�/0�d�V�G�gǕ�N��6Ɓ<V�}���p�,^�f��YM���Xcw�ga�Ի�=::t1Ci�j�y�cRX>:5զ�G����<�Hu���T	'D��8W�|sr$�Ư��bS$y"�P2���V,����f4<fG=�H
��-��m���T(ۄ݂#�����
K:ĚG<=g�'�V��a�6���� �F�s_x�['�wI�}m�8?�2^�+>`
��]�5t0嚖��sp ��_����%�q���j��N}�]O����0@o�h*,�9m^+�aA^��Gs'�� o߀�c�ܛ/\?Fȇ��o>YvZH������?��D��Z�����+ ��ڴ��BERI4�xP�)+�tù�9/���U�K����&�6ݭ3��d`݀E-?�@H�k�"������ةkiF�b�+��"�Q'�랞�=����d�[�(�[��U\�kT�ho?�}��}6�x�Q���?L��@���%aͿIMj}���p�����43.L��C�����>�h�-���RL'�i�����T�MӼ{�z]³E��5�v��2*
��@�)@̒��[X���֏�'y�F8�T��<8��=�)����hp�I��7
��]{n7�N�2�䊠#�`�bՇ|�,�5�k��lf�\���9�ۖ�sc=?��$-e4�H��e{����e6_
vj).��Df;�r:66�fo�lo��QtwEo�>���Gp	ƚ�i<���	�nEc[� ��a���S����7ÒKTE��xv�eَ�Z��
-�w�y���(���Lo�PZ�5�`����ɒ��%�-�#������-���c����J�d�'G������T`T��>o�u��I�Y�/?)cb��B;�VN�n���^��%=.�=�TC�����u�Bc
�w�D�.�������t	*A��PR��(=�;;M3�M��
����iV<x�߻���Y���	+�{,��2�϶���;l��k�.T�*��C/�tf2����8��[��GY�X��<rN�[�V �t�6�d4$xs�.�ݱs�\�85��м��DlĜ-X��ku��Ңb,}р����+�1���/O�����X^�M˗��}������~%U"�����8��!����[b��b�7w�ĐP�h�ƸNw����,sk���ak��s�-w����du1hg	0�$��)&En��W���Y�����]K�VaP��2�YЋ#�UL��<��l�p�O1��[���^�?Tpa�iRqHE���4+{���߇�]ad��]��O�����(0Eg��� �ws��?��H6��Ec�K���J�����p��.����.]��bq��e���w��X���{��b�
��S@Z�.r�o�n��m 8y�/ɍ?C�/ ����l*Bh��u�5�Sv����?/:GE$a���� ���JhT#,��]IQ�;�G���������-'U�`���c��PCׅ���d�'��/AF�
Y�F��\�q�3��v^�ӏ (g�
����^�zjR|{�Ý;=E��:=-~=�6�[6r�X�
�aAᩞ�t�;`K �G��g��*
�������n���ŏ��3��!-H�y.ͭ�\[:&���1�6����w�ӹٜɞbF���[�E��|��>1��g��5�L��Z�0��Gj&�4�P�N@�_Ϳ��?�s	�5�!����|�Zʳ��	G���O��Fv  f���R�^JII�u�V|�,�>,��������ʭ�u�A��LW����A��h)���?�}���ݗ;�N�����"\EY�����2�O��4Â�jT��$̑%_H���Ę+FK�o,����wqq�h�.�5GU��~�|�m��S��/�w���n苙L��~�?�ﵢ_�cX����j�`�#�S!�yE�#��1�>Ăn�h��U�ww����u��π[�r*�"�շ�a�]&�"�����Y������e�������o�
 =����Xה5XR\�h/��
'���: �R~�q����A3�D�L=וX�T
���_u6�N/�r�zޗ�q`� �yay%��)4��yHfN��+��"��n�$�jTѥ��M���4d����D�����2����n�l�6�>]��s� %
W�)-��w&����;g��ՍE�a�H��BP_/_�� )k� �n����������/SB`|�ܩF�R�1bDy�ݿ�鮫�o@�>˴�J�HW7�t�R��g���)���pv���^&IQ�J����̛�0���++W�֞=���T��YEĨ�8�P��٬s&Y�x%;� <��/\�1fk2�h>�ȹ�;S��*�>�:��~n�~nD���c�����*b�5�U�V\G���b�j��|�y�`fn^����J�y��aO��]��D�'�ݦ���(u���)0�
�F{��bf���\���D����R���K [�b��K��h�#��k�5Co��s����������؂�v�-^9̉����	����8���d/&��i��D	��Zc�;:hTvq)�`B���ue�����65�N�-�j���OƉ5)]޻��?���ij�'X4��'��F��a�����;C��w/�Rb���/G���>�ҳ����_1s^y=��9�ȁ�+��d�C8���qFs���h%����_Q����������4�6�<� E�@��K�ZOVc�̏R1����NRY�b^l8�H2f�Q� �fB�v�E0�]����F���G�	41Μ�*��~ z���{$i�y��Ɲ1E0�g�D�x�u
.+�IY@�rd��ځ�����gX��"��%+�Н9�ҍ��rr\i����(��kZ���p2z{��h�=X�$ɀ��[\��D�B�<<F4Y�b��r�P	��1v�6v�kLJ
����_䤝�M%�=P���cYN6��[3맅 SoB�-��8$d��6�����UQ�o��+i�GH�2 
���%2��e5i6�S�����[O�z�IQ��-��������F������Æ���y>$�Yc=��c�;��;d�tH��C��],OvI���~+�.o�`h
uE���4�'á,4���X����S�爋�ѷ�� /�F 0G���3�u��^|y㏠V�Y�Oi��4c�H)k�9^�;��|�͊�`f�- H6�RH��W� ��E�\��M��`|n��K��ɺ�?�I�5��O;�Dq�g��_[+{�P�54�l�}��ŵ5����mѶ�q		~$�*@�wV�!��j�!+�~��Ѱ�|v�6C'܆�����p�2CG��J�4Ao�ƽ-&�kƸ���u�?�)��w� �V�8�;s�n�#����@��M���ٕ�u@����#��i;w�,�&�ob�f�����$!��M�(V���֨)�j�ȥ{r��b�b�vh����ѫ��v�5�*��c�c  TA��L��Uű����"gZ��1^�/����ƣI���%C��<ͮ�ʏ����E���S5����B򅞙z��͇_�!w`��b�#�4y����B��AAAԨ'����9�f^:��@���h���_qS�Z�[�1N�1�AB�Qh���)=��
��W�}�Ġ������F������2胎ֻX!j 	�>�D��ִvW�e;���s�Fr���#p=Iʹ��X���߹w�0��ޗǩ���w���t����L͑UG\̦�����Ȫu�#@ʘ���`�:�
/�jnf&R�����ո�{����v�f9IP�Bө:�4s��]��z8��
,WA �[.|����diV���"�xkt�s�u� ���i�k8���ze�:	]/�(�K]Ĺ!��p�zna�Y<�ӌ�1A ��B���/�o311ѕ��
��ɿ�]8=� �w��c2HH�4�� ��}�A��Z�%,���:s�(�Ȋǭ����f��	�ˬ�]6x�h�����P@�J�h�g�1 �����.��$�HU���߯�����,8�����\V;9�͇�j@Q�0���BT��w���D�.Rq�lj(R��4��������p��{ ����k�����D�
:�96����#���&J2�4ﶶ��7*`��i>9�(�s�)`�&q&�r��+z5n�Z�n���o.�������=�kb��ps�&q8�W�8�����x�(�Bȭ��]�����U"R���;@�|G�ʇm���T���Xh8����U�!�X"�a�'%q�7��G�{�������s3-�C�Nz�����VJ'�����~�,emG���@*!A�ZE۬=F�LXqN:�Y��c!2HOD��c�&k��	������*��e����.>���	M,�G���+�fU��C��M]�j�N�>e��_�͉��0o��n�0ֈ2�ѥ��v�D�w^��؁�`��ڴl��z�SÔ1��.�4SS���ڬ��>�X�GK��@�ڵ��#>2����@�t�X��) > �m^]�����$�L�q� ;^?Sϸ��&�hk��bx���8�v�\�����	=��$ʋ�>�d8����$�R�FRJ.	|�a�:�ũ��:ߓb5��<�o�ϐ��@9���@�T�C�)��v�I�?r��7�9�{�m�sㅅ$��{��z�"�&Y�\E����_����G�N��Z��L�߹�tUq�#Mjj^�2�C�Ejr؜��.��zk��:�eO�MC4(���͟i
@̄bRq�&�.���&X�F���ن�q�xX4��g�#��bf�t���.֑7Z�)�쓔iɃ��Q%���saL� )b�^SPdl��4��U���
Lҏ��;�gW���W;k��]��C��f-5�R�Mox�ڪ*^�lsް��";b���ܢ�B�n�������*^�o@p����k�LP��^%%%R��>j�v`��&hR�CM�qE˹pP��4����2�ۚdj��E~*EjZ&14��Yg3������%oT�kIi-[�y��
�|������ϋ(���))$��E�ԧ��c_t	C?f��9���$Ji�&E/)Q
㻓�O���Xl�{a�ʹ +"I?V@������&�N4�|�O�.�A��@ ���IrR����D�^꤂A*� ���(^��T~X�|#D��:��L��rD�U%�`[)�$�0g�諽<R�a��`��M�������mF=���r;Ek*;�:ͦ9IBԀ$2=$���Ø��ν'�P�X�<}�zIp	��$��0��S7qyψ
�~�
��D� ���}XՈ�G���Z��{a�'��fVV~��НY�����(��e|M�nx�.t;��)X���@6�v���9K�Hp�J�{����J�U�:Ds���(/��̣�	w�o�־3�QThYm����GMR��#���Qdm��;	$�s���_(X�z�X3��dz[0B��Dm7���Q��H��}^��,P��od��"F�{�5C��@$C�(ap�}I� W�vJ�U��&�} �ۜe+c�7��P �H���Z��h\�1s�N��5�f����朱&r��/��*��Q]��JL��/~�>A��̇1 ����@w=;���$����a��:H�gz�P��߇Z���,�*�$+�ڈմ���)6,������D��O��'*v���A��N0�w��׺_� �K�`5�*-ޯ��o��l$כ�.���=��
U".}���}ٲeT�a8TUM}e����̮$�h�`D������;�UЉ��Ō>eZF-tl��G��OG5ͽ����.0>�z�J�#4��T��������1.6�K�Q'���a#O��ы�����tĳJLL����ğ/�K�sz� � ��}��M�v�����vf]��*yg�����1}�t��Km�<�(��A\��F��,-�H2���>}:�]�"���L{�ɾ�?���忘Qn�Ҹ��NH�Y���,�U��t�-����*5�E8��vw�:�?$�`�-+�DQ�B�⊁�!I�\��$�>�n�tޢīV�AT.$}�����??�|y}�`Ѩ NC���)�I%{��m�	�U{{8l K���o� .���b�G|�/vZPU�+&}�		��?��m%]K�9L�~R�b��� ���R�X�O����dT'�}��bi�+7������$��X�^H�Xk�,��H��R�V���M����������L�ъ�0,���^��U`J5����FL��R��Q�a=��N?���N�oO!0��� ����-@pr&}6Q�#vӣ�x`$uv�)k0���� Zؖd��d�H�<���ݔ@��Lğp-J/��B~;aR�q����+���I�oٜl��g�ja����ߔ���Gн�>qi�M}6$�?�;�Zj��1��\Q��k�9 �/I9s��&U�+�coM�fh��^d��Dl�����f��ڍi�g�4�E�4w��F0�����Ԍ_��T���L��8C�M2.˃FB�}�}����gb�ňTa1x����������5w�EH��R����\⴩��~'�Ay��Wz�&�d?Au�����ƴ�xP�x��:��iJ���������X��JJT6�F�fn%��/���؈�t�4�~|,\����ǊL���Γ�P��?��c�Y��5���;bb��s/����?]x9��_�:ijw�X�_�5_�d���>w+x��Hf�5B.!@�ҿ0[�d�
�ӓW�,�+�<�]�p�%(��;�f=)��~ɫ��`��/�Sy�ޯ �aA8�7IM�n	a��0�k�^]a�T�J��#��D@�	n�ձ8�G늆��NR�.#���,q�r\ϭ�s�";O���� ��k&��N�����a�+��,�d��e�Iu�qS�?���ڀ��Ɇ���g���%� �T�`�!�T.�:�n� l�4�-��е�
��OO�t�)�<��ĊV�Bq���F��f݉YDL��痗0s�ki�Ϡ��y9�8�`�6��no��|r����c'ô�n��u�q��2�eZ�H]��k���N���8��Zj�H��Aatd�*��;@���5�V����I^^+���R�{�	�Q�bt���Q	�V��� V����V������ټ������k+���������b�6������a���AT��LUTBBB�c�pq�4���%�J�T?<ʸ�B�+
A���k����$ \��o���:���0Y�?�1[Lv]��cݭ �q���A� �aʝ��0�@RaR��1IA�"��NX߇�0X3;��I׿�0f�5	�ϓ��%�	~���c��T�NY�c/�C���W��N�Ǯ@SW�����)O�h��hc�j)�=��Eʽ����z���6�Kk�T�|||�x�-K��+1</@.!�h:	�JCJU�"��E�f�� �8��m���40Q��7!���1��S�ͯo�cҔ<y���]M��U��Yk[*O.�~����m�M�Ci�&9��$b��xGK�2�B$%%�B�� �r:�(�� �3z_�eJ��yI�|�M�C���������m��L�Qe�6�Y%�i�&p�@�N�LP��V��)�)g��"J(��666�p����^	��YY�nkJ���
}x��%�n��C_�[3�jk�a������134}�?w�	ӝ�Į�n`����`�ПEC�<��gB������x:I�F�)%��Y8_Q�@:i�tŰ�����|.3��9�8��̙��A��NI���C�-�gε����4��r>��y������l,��w41}�7X�4�܄Gp�k����]�[�"�W`tj���!([A�
�(�������!DXwjCp��J;bF
�`�l��8�9����%��XW���^@���\0�!��߮�o�œZ��:����с�o�oT�w���a�A��ra��𾎩ƑA�
�D���9��3mjS�=��ȿ��%�⽚>>~?KP��31�mn�����Q N���4����t�Lue�﫱	92��*1c��/�k-'�}~��_1ƴt��-x���ԛO�?D��&8�O���}�<���wfH]�6x6�I���Ys�y���?�9�e�w��9�Al��
�~�2}ss=}'�%�U8?7{)�A��)�PM�I�,3|e{^�R��*�=�!�vG� d`��^�cv�J��G��5@������88��rAGڗck�z��;%77�ٲV�,^�`t�gA[��;�Fp�`�A7b����&�;U�8��Q%��+�y^"�T|�@ Չ��7/�Boo�I|��G|f�F�i)/>�Z/��FyѢ//�V�Jje��'����\����s�7��n�1�4�h�x�}xo�m�GS��N5���s�(�߼?kWj���_Υ��K��V���������{0;tމ-d�VMM�D����2a_o֦FDl��VR~��a�
��'JH���	_p�����X>�TZ s�.��j�����/@���.~��̋�7(ʌ!�0;�]0��Q�J%�F-�	l�r��O'��GGDDD�����׬�i^F��Y��kD�6���c�J��M�U����-�� �[-�l���~�%�s�a�wL^�C_�u�l=�R�ǡ'U�L��\-%%�uS��]^���گDj��o��/���vy��x�̦����ێ 򳅮�d�LO���?����?�f�Ut����"`A7�ď&��	P�FW�U�PA��FԦDGG_ś@D4���&8-��"3/������Ǥ�~C������VWWk28�w�Ύ�)N�!l���]
!~ڱ��aW��F��	�ˀ�&c4;D�D���r���: ���%�����fj���W=�]�f>���NJ&D�AQ����R��F	��nJ|�:wơ����������1Sz�\|i����Ҥ���ZX��ط������kl���7�䝊4�f��x���m�Dh���t��p4>��tl`һ�­�`���*��g��	����oa[�;b
Fi���;�؁�����}7H�f���=747�9�0ݮ/�x6ô����1�Th��76�X�8�Gs��W�7�F�Op�wE|�o�x'SL�
�Q�Gk����S͂�%l����L׏�H���+;L�XfƝ�����v��3�}��捕?b����w�����=uJ�~A��@���_9H��&��J<A�27�J~���ÞaA����`~�4y�3/`N�`��X5��s�wK�hs�H'���{�K��-[���Q��x��R;t�X95��;
�U2>�֌�H�
#�ќ�1��������ӛO:�wjm<�W�/}���}�zL�jE���@���mX�/õ�]� ��k0����O�'���~�8�!�_s�Q���,��<¢��A7��Iw�����Ԫ[r'�-�ކ(���*��}�� ���Z�:A���+�u��d��J$ɽ
!j�C��f�j���� 4��E�{��{���-�L�I/��DV�)ǒ�YS��z]��̭�����ӯ���ZB_"#�n�AaV�>�}H;��ЧJT�����1�a{>���������7���|Wt;�%�7���2���&ø��%f���Xd��7�`nU�3/�m��`Gg>=��Z8G~{�����8��5&�FQ+!��;�ϙ"��� ���#�bW���r2��Z��}Eh]��paz�#e�7"D�2�/HaR�C��D����xx<i��iџ�B~�HK?2o���/鉝Ɨ\���L�An<A10��0;^�*�DM�����c��z��_�zj���??a��X�j�偣>h&�f��t(����;�
��������c��=���K���?�`Dn���J�z3oTY�sM�qU��7c�����#���x�{<��������~/E��<�y�a��2�ߌ!���덄�ob�>�<��Q�^��<C2��Uy�&'Km6Ⱥ+�{���0������L���;�v=��<�g��������X��i�) ����,�ۆ�}���Bǰ�w=�Q�֫��L�?�1���$#}�\l�����������%�F���-Rъ�JFK�_[�hjy�nJ?mFY�|i^��g��1y+�m>Ǝoզ��LbQ'tT���9�p�|�ҥ�U�zv(HW�L��ȧjA2R'K������C�ŗ���=E�s?�!�L��ʑ,�ڳ:$a� zh2�/��̴����񫊊Jo�=p>�=���Te��s�pz�un=�~<P���&f ���>VF!$�0��Rt=۪|d��Y�vu��N|^����!�d�ôq��K�k������0r�r�U�����ʹ(z(��+����cl�lB��=�C�VHS��l\��n�Up
N�+�
;�V�L���o�	5����"�p��X�4���$�	�tU������8�7��/�����t^�G$����~9�N�'e��o��-5��WTTDm��p��"K"���+�m�8�8.�7�\�U�*B�41a�`�?��1o�<|�Bd���O��U�8l���
a���TЭ�yn���+���g��k_�R���*
���[w��zKuM%��w�pRY��p����ş���3{��b���Q�ZB��X�w�]�g���p.����
ȫ�OS��k)u�o���cN�ܒ������������W"`���= 2$EhBj��~�} �����CRR�H�
��Yqm��`~Z�W�Wo��	C���w_�	�LLZ���`���1����mƃ���'i���Z^�k^b�ׯ��6���OL��?2yȄD��KKz�LA�
�P�7<<m+z~�/cw���p�^|iJ{0n53zeS��UR$1[�7�Y�p�]=�cP�����h$)Ju�L�}�7����L�p�ߴ�=��V9��_۷��ֶ���&���NL���,!i���D��Lw6GG+�p�5H|�8���qG�6�rN��	jf��Joo0�O�>}�Qp ��ŇA�q�z�"P��a|�)�w�������z�H�0�b �7-gWH[� I���]64̰��3��z,g������K!V?�� l|�~�ky��P���٨i�t=a�;�U+���o��n�pd~z�!ز�>|ϵ#����3��&�L���Ejd�zR��TYY��9©u�X�ZVV�`�n{o�ZP�8�鱎�j��*�OE� �l,��p'��D���5@�}��+f6kFrU�띊3͊�-� \�.N�[%����5S�%���QaM#5V~��H��!B)�8�&��C���=Ht~́�WQ�V�፫���mx%�/A/X�@3���^[�g3o����@��PaY�������in�I�	�
j�cυ1��E�]�a�6???I3�Y��'))��5Vo�k&��F?s���"��/?�j2�SWV^�)q��_A���LK}/_�l8nk��U/e�oƨ�.I�|��v
}����UO��=z3�-8 (//U��E�d]�o�m[h��ۺ�W����E�����1!��6�9���.��E*Ʉ���|�i��O���5fziֿ�+
�z�h�u'�>%"�� ��B`4��+�������7�B��#��>�ٷA��B��=~3�|�զ�m4_,!�&��t��Gz8f]�M��׊u�5q���I�?�G�~ML�/f�\�~aYe劺�:�6nw�:��Dp�W�N�(m�\�]�����ש�О�ύ(l�ٝ�ĕ����X��s#�FF"T(z�������U!�� V��oEEH~�R�k�W�Z����N�M�S��f0�l@�wv^���i���ъT՟}����'<�V��Y���a����A��qw�w��L���i�'�|i/����D��(ni���vM�q�`t��%a4T��-_���9�%�K@��V��ǿ�BJ� ��ޓ���z3��@��ں�>#u��{����#�˛]^�|{w��DȞ��}��$>�$��FS�_��*Jݪߕ;7.=��a�acQ�!��e��N��V��J�d���_����E�~{�P6�HĪ�
]�EL�����}�B��$aQ����d�����\�(��}��gO8�`�pҹJssw"�,S�TQ!�׳�s�A�"��>ԇ�ǎ[{���I�+��5�-�K�Q���`g�`ׁ7p*�d�*�sڂPD2�љ���"�3������[�� ����*���ӕe�?��bs�ͧ��6���7�h\�������=���_Ǚ
v��Y�eL0��zV
��鞘U-�ĩ���v ݧ-Ÿ���3�k�㏽9����jD��<���@c��{�_:��Gl䩛��Ӝ���$��0NN�+��!�B���eT�'臏�c_2�O�Q4����Rs�_a�c�E���l�O~,��Ϝ��w⌋�#5�����Ok֮�{'���f��짮U�ߴ���r��l8���Y_�|�,���i>uqA��#�,��X!�f�:J��WPQ@<g��ʨ��Y���~!�!L��ǀ�B[��P6x={���T�6����(;g��6�Ź	�ш)P�Pc��?D}��j	�%#0bg|�wͅ$#���p�(㙄����P�aأ;��,�|�'�<פ*�ƘP��؝��M�qףd@]�/��[��2?5������I	/�:���A"A�H ���`a~
�\���.F�L�<��ŅL���Z�փ$i�&cpmP�U�`ۋ����q{e�*p��6�������ͽ���}[�SӢf��Gd7��T�2"�s��bY��)�w*�������ǻw���qI"����^o�)FP�ŋN_#��V[�!do��$�.���Y�1\����I�����an�����Ltx�|���!߂9ɕ�X��Sya�B0-��`���=�����G�y��%�.&rc�� 5�����SV�"=ommeNK��@j�����h-���֟w!e��Z!�"V]�Bd�m�vV�wuyc>n��a�K~x�ٴ�`� ,��[Lv�D=^�wW'��Y��	�*�ӹA��i� �ga!ݰb�%t���iҴ���foX���>4�"K�_I����c����>��a�t�����hT	�>��_)*��o}}=���@j�-��A���
~�)�����r�T�,e��ѽ��E�'6�!�~o�k�yl�`łL,Ȳsp�(�!�����/������xˇO��#+�Y�h�b���`*z�u����$2�ϔc@��0�˰Ot�Ǐ⨣D�{��F����0�@%uw�~���EI��h������u��={��̿'a:'H�Ѽ0̋[� M ��T94_�8�X?u���pU���o$:���3�X��������ZB?��,�?^�!��U�W{�#�<E)�һ6��AR��������b�4C���z�j�����}q8��`���à4�0��9-�ĵ��x,��H
�nC7�%��Z�<���L�ʆ�.ED��	�Z�ti޳R��LUgN�Ɲ�;���D�:uꯠ]Y#է1��.��1H%?6.������_-�����F�+��ԘFVYE���J٧O���rPA�-���x(0�P`����1��ѱ�P<SL�����
ڶ�� 
����`����Qc�8&������B�ۀ6	j�H���Y�;L�`6�2�;�G�ӱl��L�cӈO��g�����rr���@��J������ѩ�Q2ߛEm���)ժ!�5����@$w�L@\!�q�o����]��򮇿$�L�c-���0��;����wj���Ԭ�d����*!:������Bh�c�����R��̦;��o��ݰ���;���k���RS��?�*U��x�Ԃ��Ʈr
�)�,��1&�����28�ڷ��'�� ��7�R�0|�]�r�����&?�(�t�6{5>�f8:���^*���K[I�5 'O8�|��u�믉�%y���24]�<�(��3�u� ����� ���k1��ly*s�/���G꺈��q��s�����q֧�OY��>e}��������)vU'�_r�xt�u	����;˃�b�X�����mb��w���j�Z���j�Z���j�Z���j�Ok�}���q]5c%*9b�?߇�X-V��b�X-V��b�X-V��b�X-V��b����2�����o3/V��b�~�t؈���y��׺o�x��X-V��b�X-V��b�X-V��b�X-V��b�X-V�rk�C7yL��uڰ���5���8Y-V��b�X-V��b�X-V��
����w� �m��j�Z���j�Z����J<]HЉ/N�E&�m����+�;~�)��j�Z���j�Z���j�Z���j�Z���j��lї������~_½5��Ĺ�������c.Z��׿.����;��)jm������������������b��5�����>~��?|��Y�d��5 k@ր�Y�d��5����kzz���م��5��*�ږ�Kt|��k��<�f?��+ެ���!��.N��]k����94���[}�缸(�ߒ�����������Xqa卤���lO�iK�y�+)Ŕ�Y�+gP�}z���g�{���I:�mZ02�E����u�.��f%ۧ�E�GJ��&KO�5~�a��I����O��Jac�0�۞�O�^F򎰓Om�έ�GW��|v~.s��ۤ0���r��&!8��z��:���-EI����coO��9���c�.r�8E�����e�ů?Q-��x9�����E�F�=��>s��&^"�����cs�������:�\�����l��u���x�H[k��F�f�V/N؋VT�z����1��_���X�7��0/�͉3=חYԴ�2���D��X�����j�������lΪ<X��8r����6_��r戡ai��O��ZTӂ�lmm_�)��w��,�z��tS�y.����̝��q�ec�=OՌ�o��>?�����N|�t�����%��$�a:�t��ٸy��~����>7�_���HW7�k�� M�;ǂg;>�R�Т��7�ו��46����̭8y�^�/�%i�Iod�@~�-�W��E�5nc�M��$o�Rt+�u�l��i�A����jV��:g�K|9V$�m��� R?~l�L�.��/��;�� �o���F�;g6��-�ӧ�'>~�������
�m��)�[��L�2�~�&==]&\�A���'=!>�U���Gt���yڸ�٣�����׀p���Όq��J#:3�;���ڿ}!,�f�y�\'�VK?����t>�a��3�ڕ��W�mH�5��[J��Ţ���O~�ٕ�
[��G�pv
�	�͖z�t���$�ky������b��}ʀ�{��v�G:�6���_��^�{�d��B��7)�m^����f?E����k)�ms<�olf&R�(��I7۫�*��x]m|H����N�뺉6����]/^��Ñ��Φ���،tU�Kv������K�����2��.J�x������	�T�Ġf_�G�^�G�3�}ԙq�������\ⴹE��k��+3kA�]/�P�V��Z����@��>����^J�nW�|���xk�ۄ�YSa7�>}S+9+�E=7#�]��	U?�[��;�u�6��{�+2��c^����;�-řF��11��H��;��J��QHk^���3#ͩ�Hn�=̦�6���nq�|F��p
͵�6C_��9֥ɇW�t��ON���4�O�q��N����}��6����@S�j:v�����+��efw�E�B�#l-�Ͼt	F�i?M�����fI8�kz������4ڞ����NjKuixCo!t�����ʫ�Gw9$�e�?��Q���o�Ro�dKB&��o�O�N�iJ���q��)zy�O�>m�y��ѫ�=,��,}��k���V���A�Ӎ��w�5���� ���କ��=fݍ��sMlF|s�-1��T�6ǒ��.�9��!��_Djɒ%�[����t�4Z�^�8��у**ð��IfJ��;zG'���
>b�O�n}zbRүbbbt{��c�k��-GYK4,����N�h������`[�Ao�#a#777zNK�e�ԇ�6_?��;'Z5�|J�2�1�jp�2F8���Mv8�^ͻZ�k/Gyy���	w���������Gdm,��T|#1���mw��}��;&��{�;̓��T@֯2�%''��p�wg_,
1��IIK{�x#�������Z%SSS��Zm�jj�������V���ݹȴZZZ0�����t̳_$��d��d�}a���Z���=���L+�k��G���?�`r4G�� ��ɑ�k��çj�)���4!�6g����F��2������8{5�󄄄��`���c���읾5�ւ/\�~hܓ����C��D|S���O��*�}��mm>4�T�L�>yy~��V�ϴ���oLA}KS��IB��o��j��WY�h��t��u@'��`�l�!ضQAQqv,ѸP���pL,M4&ԧ_����w�;�LL�>|xmӁ���4��/���6iUf�ո/ق/�L�U��_�:�[Z�,��u��o٧j����S
���1j�qۺ��Y�&��e�5�i� �<i�q���w��i�O��b��;�C�u��I��*�>*y>]k2�u�BBf��_}nx�lYm[[��sק�%��n��O���+�׺�u�#�`�wZ��y$����kv�f��#_36wd���I�ګOO�A��m�l���	ǵ/5��'w�^ �P�J_ۤO���)����͈�^AW�K�b&G?.&�g����C��S���x�Og��K��<���C�}��˫���W�g�ߢ��i��>�笞>}6I�k��t���>�L�������'���t�G�11��\h5>Y���m:��^%�c�jI{��:�[%&�2���c��;�7P�w���i�3�:~��#bbr���{
bm'�sN��q�
l-��ˑ8�86�Sth	�s]�p.�������e��b^F��}�˛��5�<	��Z%[�P�����G�6��}���c��=��r�Z�M�Kݥ@Z����-��
F<I�*�5�'�j���0[	�I��I��0���t+L��=��w���q{�/<�Y�jn��I������P�\��g��ٔ�ՠ�穕kV��r�2{����I�^�,�֞n��F�[��3�E�t5�Z�ͼ���N��/>�{t
�J�)����Ŷ��������I��2��O�4����Z�Lw�I_�*��76f�;�:�a��(�zy[��#T�g��~�v���h,��S�V��{ԇ�N>�7Շf���wG�Z�r��_cl��,CD�#��	�F���5���(\|v0o$�#aw�bq �.��!ɛ���tw�O���m0���E���������ޙ�gާtG���+V��EŖ�rӲ
��ތ����:��=5���d�nS��&]5�V���j�=�9p�[�-�� ��vg�x�4���ڷ�@iK	}�߱x��d/�#�3��ʄ�l���"�C��Go��JKJJ6����4�s�5������XT�����bZ,RŜ��=u���+��G>�~ASfC� Z��ԔU���8�9�~�T`+�Z�B��L����RP�ڕ�J{��N3�e<0bG�ӧ}��̒փ�'���"�B1k��Տ���#����&�<5�q~}z�e�0s^w��������&ؖs)g�;*��3�g��3��M�}];�ӳ)h�䞨N���>ڻ�%,bn�pB�"�Bސ͈�ğ����tv�ff%�)*�g%[�m_�#D�M���i�Spnɽ0/zc1�j8y�XV	O�X|�<RͰ��v0�(s�+��C���5�n������ӛb���%�ҵGN����s��@`��-�0l���ƭ�%R*����g�t�C��D&����m�>�e��צ�2�&6u��W��O��.�4|���qd���>�6�~7��\�S�3����Z�"�����|���ۧJ��hv穔<�1�?o��$�:�ڹ����4
�x���7G��i&��g��ݛtɮϖ=��=E�;���05��@6�K�E���RD�q6۲c� ��Y:���R�w�?���t����8k׭=y���᣷#�������G�f�R�j~���H���HM�R{�ܾ�,}�cǜ��c��}-�iv�q����ܻD���u��n=��uqo�^���)~vN(�b.-w��rI+��Wzߑ���3�x���k
��͢u.��!��^v�ҥK��@����ގ����T��}=�I�#�;'F}j~����?��y7(�m�ל��_k71���/l!���wH�]��լ�<=���	�GT���~���#G�d	)e�nDRb�z��j�H�w?�.�l�I���l?��m�[���I�=Rк�"�F&3�u\Nh ���'`�U�/0ia�����h�mi�#�z=�K7�6h�r�$ׇy��uh {�}�gdZ��^fg|f������L��������Sͭ�v�I���p�Z{����vC@�O�vdXrqH �ؒN
`:���5�96ԉ����2�ҮN��]688(Dּ�{<W~mSW�3׶ Ǐ`�߷MeΦk�EM|��l�ӧ�rH���A�lܴi��yĊT8>3���m-j*�N�4�yl#_Tn0�_KQѺ1����X�#a�h��5)j+��{�Њ����8��B�����QP��{��ro�����0���x�&�N%���,�	mN�8�m77�Y.�a����/7�>���Y�V��^�#�[,�}PpT��6��;�?�U��6��bY3{?b��o�Y�(�����Wi @�q�Y�,��m83p�þ\���^z�;D.e��*��rX{��ޞ�qg�����}��:�~\ץ�w�����-�)�-|uv�[@��\z\��=L&��N�Љ��p�`L�m�1���g�,��mrt��og�8�,G�v�C��ԏ����P�:�d�J���ه��0m+�z}�]E&��@8��-a�������W�tF�k�񖜣�v����g�� * Cq��h�#Ge�^��-��Ϯ!+=��P�U`P�<� P��y��-���v��(V-H&9��xl�Uԉ]]ghf����.h�;w<�`oГ-&��q���I���n�n����壷�{����	.y:M�}�����mHWϞ=7�i���P�Fi%7w�2��7&/î8�h�<�S~9�)���q׮]�N~��=����WWz����b:�~�:~�*t���ם&���2X0M1|��X�x����L�r]�&�Ӣf���˗V-��o�s~���Gh|�nP[���S�� #�U�uNՂ��ګ*F��N�w�0O����s39��,ԙ����\���^�=o��YM�`��d��:��w���#��i ��Ig%�=�+�	L�՘:�@ϔwd�ݧ�����:��E��&}D��':����6�17�-U��)�5ܰ�w��=�Ik��:�+��}����������4��֮mAR�^Г����:+��ڈsv�7�lG5���s8��ҲG�G x������CJ�1�I{�-�;2#^4V�j���B��%�nKV+������~P���W�ק[-�T�Y���wc�}̫+�L�Xԏޞ�����N�r=��{�����{�b��6�Ӌ�a��:0��G���.�B���엫�B�Adk4yӬ�/.d_>1=� ��Zq��/s���O��TVL��	!�pPf�h���]����v��7r���P�tn�ZH8�k����w[�;+�u��-�6+@�uD@!�G�*��[�K�>���T<�#D�q���'�g�߾{��,�\K��ಮ�.��x5�u���ޚS�cgA� 3ܴ�|E���8rğ����>7�����0'���m}zĴY�RG��=!�i2��Q��I��;.��M���z���ɲ.{kRN[Ը?�wf�]$t��:�� �����vefL̄)��~�4�Kwdl;Ƣ����(�s�:��
�6L8��?��q�Omm��sC��,��w�c{�/$ކ_5��ޖ�)5pq(��rF[�b�<�!D�!*��fE��A0+�E�����ή��0+��5���ka~h��bX�������e�`��l��+?do�9(QQ��n�����q�Ӟ��ys�9�6|2!�k[����)s�ɷ��S�n��W���]��OI�yl���M��ʙ����e�v�M����v�����y"�o�)о�J`z�~�+��E�ne�k�Lм�)�v�����b��3?��3��"ϝ�3n޼iL�^/ϦF�[�j��"sh�>���.����wM�\z?:2�����~k��&Єג;�������	���8P�������i�b�6O�^{{�� ��S.����ۧ���N,�?��i��D��4���v��?ƺ�٥sz?0j�-���r�~�����]�~wO��~k��|u�y*���>m�zfkZU_9m}_�z�ӟ\S#���}�L�uS`��C��K����t
�O���+'>8�[}��B����}4�F���^�c09�EN�ܪ|ߖ�{䕹��.u�G���I���{��3�%6�w�Kk9�T���^_���������{:��������^<=|�4]���ze��iͥŮ�5�K��ܖ+����~��݋�A��N�;'��ʾ�ǖoy�k��)qB���S�
~\�H#�_�n���}3�No�������}U�+-qu᪟u���]�����c��9���e��ү���z]I?W^���d�9`�;�H��v��f`�ڟ���J���?�_�SjYn)�(OW?�uN	M PK   �i�X�|�	  	  /   images/e1d4e862-170d-4bac-8b1a-e4319ef50e6b.png	���PNG

   IHDR   d   "   ��|%   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��h���O���&���1�T��]W6�GeJS
ҹtD���m�f���]�1��R�,�9FAA+���֊�2��DI)�6m�1�5���������\�{����������s��<��y�s��4�ڵ��X,�V�X�***����U�7ܗ���<===}�֭[���4�IN�:��;IH:333.�T��l��EȬ�W�7ܗ��Yk��ּ����_Zh��Ζ��.L�B��fw#&d�t��������ķ��������q]����^8::Z%O�r��/��Ύ�q�[!��l{Y���Oݽ{w������nrr҉��۷o�&b��P.�xo�	"#<55���R/�}D$<'w�f/���)���/w����ϋ�Ú�#"�$�|�r�E�{��D��i�ؗ PT=��g��Od�ח-[�B
��v��QWW�m�"����P�c bD�a��Aqq"�/_!Me���DU������92)�E �b���3c{�{M���������P@�I�ɧ��J�$�Ab8�%]џ����ا��ғb&�u`��[��=I��E�2��8���6����K�%��=)9)�O�(s�\���>3y�Br�����2dr�w%�}mOH�,i�8���6����ԥ���\�'#������v#����F����3A���Tz��;���w�� ΃�876;�ֆm��I#\�4AEZ���<#�Νs;v�0�ޕ����ܽ-�Smȥ�J)��댓LkF�|`|�{[������\��d�o�T�CaD��{��}�H5[&���l�g�u���C�n��k�p�Q[5 �H��Q�w6v5<<�A�3*޳r�JW[[�jjj����s�@w�`�8��N��  �W�Z�}'#�?���\��ې	�T� �!9m$m�,���\�~}�ڵ�7Ƴ����_�gƓ8Dp������,��񻾾�555y�GX�����իW��h�����h�s�6x�ӏq�TV�\�J��!Ni�>�㥀+��%���U/�Ѐ��xU�'oi�9�g���LoF9�}}}��͛nӦMn۶m��ٳnpp�ف��Q����x)��[��ׯ{Ě���]��l�3�ׯ����d�|Υ���2C����;/ٲI����N@�.9"�$g�ʋ�R�]F�\
�h�L��JXB/����������$���XhCCCNi�^���$�Hd�
��� ��9ق6R���2'��e��t�Nc�#B� [NI�@�E���O��P#�-Ƽ��,�e�w���$�����®?�;4��f�o=���b�A����	[�a>[��E�2~I��YW P��Y_X��I�a�n�rq���
^^u��8k�2�S���+W�T'�6\1�
SdX9�n�800���9� ����*^:���B��7%�K�%i�fF�b����AW"Fe��G��n���8��&�@��:�gN���%���IK.��8�l߾���	wX��o���I�����EI�ZEI�J���^�ڭ]��[L1]�׳7��u��Ϊ(�@�ӭ_�>���@�=��/h����)df$�.~��?��p�����k�yCA��@������7^�q=B02��#��Bi�B�a#d\�l�<�3��Ȕ�T��C�R@?�q�C��8x��L��aez�:;;�� �&7�� ��ԟws��u��ǣ�����?n,Bh�9h��Pz���*�;v�X�z�\��b�V���#D�3�Ȑ�>r?7!��u�t�hkD������	9z����ݻw��+"8�<��8#p�ԕ��4�`6���A6j�:�Y�~j�$�{E���]!(��}��yJɰ�sV�d#[�bD��#s���W��K�X��f5��� _��hߺu�wV
"�r�Ν;��w�?�x[��UL?�Lo�SO�e�h���/o�Mm�DyUu��>��[ѨwvR�p��?~���xe4�>t��ok'&�1�g��~�Ns��5SS�YoSM�W"�*x���C����EÞ=��{���������������������������n��K}6�xT����?�&'?z���3��ӧO�{����>�ש�=)+�\����W{{�'��{V����}_R�X�YB�X"�ȰDH�a��"�!E�%B������#�    IEND�B`�PK   �l�XS�X'  S'  /   images/eb6b75ee-ffd7-462d-b06c-ecf58549be32.pngS'�؉PNG

   IHDR   d   K   �"�   	pHYs  N   N }��   tEXtSoftware www.inkscape.org��<  &�IDATx��}ip\�u���_�+��$���4I�TJ�(Y��X��Ď�ĩT%��)O��xf2��%������X^�-�lٲH��h��DQ�\���F���7߹�6Rv��ܪ&��ݷ�s�9�;˽�w &�,�$0�y3�� �cc�>{�p�g�U�V�?�b�6 �r�30�ilO$�i��;��?n>�(2�h�&4��Ɗ�}uo���L�[A����<p Y�d'�-����!���7�vM�X�޳�?�!X
�Y��P��ø�sW>�	�"T]������,j#���v�R_��-�ݯ���q롇� �7�\	�׋[�na�����?��/~.j%=On<� L���ݻ�q����<yg��0@.ɐ��fZ����Oq��ELML�c��z$��/y�k8�'��G��5��zi�l��F)7aR��
C��y�OM�|�run�֭8|�0��)r~�~ =][�%"�v���}�C7P�u��&��l���l�Mj&	ҿs'�q|#N��R��6�ӆ;]C&t>�,�}/��F?���SOa7R)5��FdHߥ�u���+��ߏXkkQe����r��� ��a�����x�"5�3g0���c	���L
)�p�g�����_W*I݆��LF�l����Lf�9>7�4B	�z�TY)�i�l-��o�tH��x�PϞ|2c�#f�www�{Θ��38G2�>���---�s��и@i���(��z.��#G��?©ӧ122�����n�F6���s~�.�X�`�"�0_������F�u�$Xi#�A��
�Q��t?����ÒW^A�O��cXEuX6�C��pS�-�q��,�?u
9�}��Wo��nY4��q����Е+j�T2Ef�(9����Qx�1XDlX+����"���ff,��2��-��=��ֵmN`ͦ�J�dR��g��״��9�v;�ׯ)Fja/�_�/�75��L)q^��؆M��UVEqrP��:#�Rp����4��Y�̥a���3K����<���QpYS���t<Y�6��}t�Z� �i��OP�Y,I�ȶ���@��'E`�5�/���$Lр������x<�b�kյ-�!2qZlS��I��g0��c�@����p��kqv�� 5�V��>�-V�,V���XBmrR���Fxj8�}|�߾�M�,S.�x�����$�<���N�S����U�X�7�v��0�T��w�!꧳S]*L&������{�����*jI;��m~G���c	żo2V�<����1D�((r�<i�g g����G�8�Q�Ot��u��{�o_��$�s��H��菘�:�8ᭃE w>�X,
��	����
9���>��
3<�{�}
$b���M**�����������q~�X�8ɐ�Yk�������c0��c�����#H%'�J�#諦Ty1�
 �>.W+�=��v8>��D��_�C&�Mg�A�=�4D=��=������w-�v�&�f"�ű�3{>�kA��(&���J ��d�y:oS4��~4-�Se	e�K5���PTU�s��,̍UX��,Ta�H�6e��`w�0���F�^Iek�O�h��+׉�'�m�&��%rQ@�vY�Q|�]�k��i-u���~	�!K�7����f1��Ů�tt�ciC-ִ8��W�`�a18,V�L����d��m_*�P��<?{~B��\,&�Z*Ú@{7�ť�+p�ul[��T�(&5�RW6��toѿI�2X�e
yW.6a=ݎ\<�������=ͱ��Wj"2�;�K�!/N 6��7�p���|��ޛp;�9L��:GD]yȐ�ZI��/��Nzَ�6ة���<O)�W�&��k8�wm� ���af��O��h��ճ8w�2�I��	�wZ�4t�+6�}���DVۭ��u�����vz�!f	��Ʉ��9i'<�(���s�Jx���eոv�U���A� R�*ò�u�� �u߳��g�_�U�*3�B[��6І�;:�9QR�}�իh�ΒV3F*���@ʴcߦ5t�����������i[���/��	![��0������'�Ee���Z�ha�7���Ѽ�޷�u�^r�<��c*c�3u�LT�>���� �t��Dج������aЭ�	��wѶ���U8�5�gdX^��=���[�	'��!j��M��@�q3��B=����	���4۱mv�؆72X��3X?I����a�K��?��~?t�D�z;:��q�P�r;��Y�F H�F�5iT�xo��+���2z-<�y�"�Ɲ�TPG8k�c�m�g�Cf7��p�Zp��\�;�!��*D��H��۷���pz}8y-�����'1�Cf���w�Ö%"x�͛��'M�P��FH����	��<��/�lJ��Ï��_%�#���_�ln�P��E+����h\�Ӵ)�G�TX�6!G�([]h9��1�7�J��͉K�'�r�%������%��|r�1*A�0Kѫةx�bW���۷�Xې>󦺙�F�`��Uah�y	�r���,�;_�������H��!a�\F�hĕ�IW�a������N5����AX]�] &���pP"~o�2�{�f�4F-Z��υ��S����q*��D��s�~-��l���ķ0˳��f˽�Z:>�N��[D�1��ܝ����x>��YE&�XS�����r������k�1���1�-�%�
b���fi-��v�N'��ۇ��ZX·���`�=mN���keF��x�fu�!�$i����t��O@�D�1+�1��cXN���ַ
��θ�{�`I(���^�&�%,�� h���D}
��Φ��+צx-�QJGC]�==x���8p�~,-�c��uE����j�=t!�8�g?�1l�;�IFp��EcND$C4�948������Du��۔R_��ɘ�uw��O����^5N�}���nN��⫠8�"�E�Ch��^��W�Q�l�̈́�v� :r�(Zy�C��Đ r
�<���Z�PT��*'A u��Ez��G�Ao�c��I�?*�(^���`�-�K-�̘e�5Mb9yD#QŬL:�U���sq�,!N*�������n���ɓH��͙�9�vcec#��6���U�`�G�w,:�t����Xn_�U�k�Q�::��Q���wh��Շ��-;�|�2� �zo��������ز:�+W�����������q_dMS�,�1	m��d=���2S�b�I�D6�=a�7�"K�'�K݅�a�
�sL"0#o��s۶lBo��汣Xu�<l�~�RU�n��B��y������jT�m����ELM���_|�[�=?�֕AtOQWzZ�[L��6XW�U2�O����2��a��N�T�G]oLL@�[U�Nd�.�S�ob��F=��D�G$$]&hc�G0T���+Q�BgOm��z�ɳg��¦��zKy�yځ4�ԩa8K������fs�����LRJz��Q�TYv�Wq?OQ5Բ��s�{V�@�"�[��z����Zh��2n�	���4��(zɣ[�������U����uN;�d�[$�k�ő<�L���՚�0(chw�jK���z��6gh��9�M�~8�	�p��)+Q���x�j�l.�;��!0q�Z����KN��\�PjB ??;��Md�)O#���T������"�
�P��[G�>��S*�h��Ҩ�sDSF,�&}9vkhٴRg�|���\���@��\��R��t�)�Iܘ��>��^����੃.7��8m��p���7hH���J6��[��SI��隦��ʐuv���yJ(|N)(��#$-_g��.\�$j��m���e��q�4O�}�]	�(-frRA�B)�!LS!�!��du����_���݅����'�r�4UV
)�kc�@�D=!X�uZ�(�QbfF�t��A��*7�.�ʁ���E�$�>�ykT 1��G�/�$�0Bc/C�+�uK�Sz��W&i
n�5�!��{�"w�&=u+���e$q�|ZZ�s���+Gz���(�U�Ĭa����p��F�U�"�;��K{n���N��*�Ec��j�!�IX�n7Xm������x:�ˑz�)M�.ܿy)::����Ǯ���8r��f[��ń���QN)��[O>��>�+����έ+�BiU
����3�+$�;��P5j��[��!_hY4�z����-[��
�!�I/|��-�vn����K���bp^�8�DT&j�����Rв]���!N�/uc,6�q�WA_]�n�^q
39;v�C�cO��6��!4	2��.�H��0�_?Gϛb66���.U$*�U|�M�Ú��n�L�u�.z�A*Ҕ��b�H��ؿ_1$�u}r����2/Y�����ӉT��T
7��EǥN����ԉN��.�z9�[��ONN�	n�U!~�׎�,d:;y������0�68=^�\.���L�HjZ���V�4e�������nс�f?ğ�d�B�r��V�%�-�)�5���5�m��M'0f�q`K;.u^& 
 
�VGJs���$SI��H&'���TQ*��J[�'�~zM;������C���>z��p	�4�����!8��aC�R�Z�0b�4HG�f���$0���b�

��?��I�@�Q�c��!/N"	V���Y�yQ�	�Ë�C?׍*��d:���	L�dB�n��l*	�ˁ�{�`�8ћ��o>�5�]�mݦ
'���A�!���N���QTQ�Z����h��>dN���S�<��`�'��}	<���@D(���-Gb�����Ni$�N5$Eo���,��(�Ef�"����OD���f�=���*H���[�DtҢw,��޸Iu��d����$n�,�Rj��R�O5���О�z�6q����ڨ�\�nRз��@�JQVƃ���1�X�*G"�%�q������ŃW���Z��wV�2\��/��V�cU%�����8%)$����j��-�9\R�KYt-�.(��(E,+#����S�Dݑ�Xb�EQ�8�1+-W++��+y��Q,s�f���;N�+�$���P��bn��gTQެ`�*�3��ѳ�M�Yj�G����8tF�&�p6O������%Awiw�$V6�K��*qy\>�+�t
�i5�u�TYv����T~~��$s����6����7��kC_�4�p��O�)}谚Y��6'0EO~ ��]V�T]���ߑۼ�LX����_���/bt�:t�?���'��C\_Z'R��JL�2�-��B�͆���i�	�X��+��b4�d����u⡭M��������%�{:��#ι��,U�.+�l7��KS�	5^�.��ի�p�t ���1�m����z?z�G�}U#")Ϟ��Bu]1Ｌ_�_�SSq��QZ2�O7Z���--�77���_[�Zũ�p��^"��~��h�����/�s�d�ɝ;����}C4d�)�[������7�;�έ�h�$�(9�y����B�v�׸g�^��Z�:��g�h���V*��?��n������*�"��R��2�rP̦eU�vh(�X<EΏ�4e�=VJ�j�
�J����B[LV�6E��)ה
�ΔT�HB��_ �ڙH�!ܖ	z��t��wf-��2G�7���n �QZR�z"Z]��B��%�+۝]W�СV��ێ�:��}�K�PU����T]�ݜ�۵[ť�J?�s�S�-��!e��x?#(��
`b�`�(-�b�L�KzW��9Mr�J=��I�zY3���ԡ2�+�Qf�Ĥ�#��,aw����`'�z���z��ۆu�kq��5�E��PCִc"��&�ʧ���!�.PW��U)�$�5��h�h��Fĕ�T,*�����K���Fb��N?��ٰ��Eu兇��I��M!�C��K-��=;������^D�X�m�EH�nP<��]�A��Gڼ
��D���]����z�d�q���):Gџ��N����RE�䖺3z�j9�k���'`_�vNFՇ�7X[�*�{������>��T]���jC�ъo��C�+�׃p����%'Oeq��<U�غt5a�7o%���/2�qiq��HO�ު4婓��x�QK��ޘ��R:pkH�:RF��G�L�,���_h:jv+-G����Ӈv�t� ���۵����9�ĭ�A˗�7�1"K�:M����`"�@2�+Ք#"���@����qX�b०k)͊�N;�qz�'O_�í�������b9�K��c����H�E&�`_6�*��Q���ȫ�ɗ�V�'����2���m�������QXsаy�:|���3���V����Nu�R�l�֍�a̶ܺ�1jmE�咷g���nɀKΜn~0�u|�,���}�zD�����x���E�½c���gc�;�Jz��������Hd!tu:�V�V�'T�Ы*�U�Z��J�U7]�����mm=`��o,6��ڊ*/J%�ni$�)���&v�	34<LD&U �IQ�m.���GlB����xz��vS*B���a������bi	R�G#�g`@��t��d��x��M��.���eː�遫΁w�&NN��N��C|�f\���_����!���.t�J$�_Y�������oK�"�vb������&U����ʢ}e-&��� ���苬]QKx�!]m8�~����LW�5a`�0��| ;=հP%�x䨪Am_�AA�rI}�w-utl�����Wc��"WX	,"���$�.H3�9^���U�v�X�⣓��舩셋�I�u��cp�xW%cU�C�ܐcW�;d�*%5(Z���1����LL"I�!�|�t--S�tYi:Ht���O��4�i﵅ӄ�WȒ >�8��WvC�ǥ��*�K���|y�J6#\�g�[�xWi�P*����*ve�j
�r^:�M��XN� ZKV��j�-��G��d��L
�.���	���Ks+�UmjD������E��͏�kנ�R����σ}p[�cXj�ʝ���(8p ��VB��.�?�i���}�3��%h��'q�����G��Oqn٢�G��������F$��D��L�34���i²��D�7<�o�ė7nİ˭$h��������Z��g��3���M���x��j͵�ϡ���N�&j����Fh*���ka��F�-V,�&����H �*>�-�iR���3��V<�?�m�$>E}u5��[���1�^4J��8����<�}��QP�!��>�汬TE���RK�wG�K�c�Em�Mi$�����Kald�+��$��2�H.B����[cz�n�˪+��"�\p��7�E-ͳ3���L��*�ߥ\��FZ����Ũoh	al<�S�����	��Z�0�����A�-����D2��#:ަ�|t�쟑�{�6�W�����A�
�\�]��.�t3�6N��'X��t������T���ʘ�;I�S>�����f�T
�������z�� L#��јRSb��x������RS�,�me��iԇc
��g&%PJ��p�b.���R�(�6]���,�lmo���ʭ2���C��K���*ҥ�ČL����N@�*Jʊ�s&��~��2T�y,��	��Ǯ��c����҉n��L����N	ɖ�Ztᴕ��(�C�8J�����r%*$֦ۢ���S�h��J�)�����C%��U��Yq���C�*ˈP��c<�������d�I^?zT]��|��߱�AF��a�6B��mG�j�J��}d��1|�(.���P��X�	�"4�����lF�[�텍��C�Q��q��^OH�o�R)\���z�,ؙB\ˢ;�D�ՂŴw��G����U���Y�ӟ����\�Lǹ�(5%vEF�����Nhts���L�����`kY���7`'�Z�����z�,
r�2Bs�V"��jm-Z���:�zzz�*�@��R[`7;�q`cW��c}k#��m�{�&
�;�n�0[Y"ʭ����l�X.�S�s�	>�����ȑ!�TDmy�Ɩ$N�9���T�"��l�9�^�l�;u
�Y[mb�)ܸѭT�n�gl�������2}�{\�s$�1��"�#��j�]ɖD�^J�������,�)!7	�jD2@��d�X�����F������Ԝ��RbD^&�<Jk�N�2ئ)k�tx�.Dcq8h�\n3�źݲQU����Jv��Qk&K�9a�A�"�2e]������+$-K�I��(��ß�ݨܵ.O�Q��{�A�?�Q-�n#0�����o������6`������A�*ĥ�g�Ù �]j�E��i,��X6�z}�x��*5W�BR�F�����gǫU݀8o�q����ð��꼱.�BEaB��ZZ`оhkO4Nd����0C�.�-�T��h`���h^�:z*g���xq�;/���H��D;��a4��߼H�شR��0�2�SV�9d_�Y��6ـ��y�ǷtH��ب}�h�����v�PQEY�f����|�x/��1����RQa��]	�4w)�`rNʌצ�
g��
��ʑ^S���8�~.Q��͐_�����q�;9�����d�X��;�PaV0C�x�y~*�� ���9iz�Y�#5T\3͐}�{�i��`������m���8�v:C+0({��������T��/�<��r��z�Y9>��e���h+�sv�തί%�ur��SL[��1U��Ԅ>���ʕ(l�;"���-%�X(G����Ϣ���%LL1M%S|�������������u�j�vЏ�pT�lA�`qY�b.�������ӻ�iS�_��l.}��H�|p��ښ����$(�m_�Z�S�z��>Ĉ6�)%�i�%�.;�?~��6��G�J/u�	���ٵ��o�PBzi��B*%����ګ����.�z��ٻ?�A�)�m$��={�� ����~ᨪ�'OB���׮��D<p��&{��߿Ͽ�"&�lA����2+�&�b���/�Ɏ��-��܂3���4c��,����!���$i�˽�˖���{8p@��*M~�B���'N`|��Cr�l�gg�iJE��`E�r��ҖT�2Yu�����W�e�ԥ����r=��ve���3��H��\S�N�&Js���(��ߟw��1�޵Q��Ґ��"1����ZXe�Y�Q���c��,V�sb�_���^��7++le7�_fF���Ԩ�V��`��d�-qq�/!K�����;���iI����~�E~;�7��EeH��J�\H�*'i|�M-�����>��	&�1Y�-T�_%!n)gl/�r�N	���N��_����o�װr���->���M�.[�V����ఔNQ]����z|�>M�رQh�t4���B�Y�ȏ�	R���N�QM�5@Q:ƛ���5J���^S��Q{�
ϗ��$QC��H��_�vc#�m��%M�:E�ӱu�Bp՜E�ˆ�]]��[~ ���{	s
|y+�E);MdȐ�W�Pd�ķ��7$�E��ѿ�[��vP����7����w��m,	�Ϝ>��Ȍ�m�Ut��"���6{�e�͐��}<~歷�$־�F1�$,�e�G�/Ǐ~�c���Ǆu�(���73U(����,w�I� O�RrQ��ƨ��$�I)�=�\�[�8�0Ml�T��d��Ee#,T�Q�\��BA�s�:�_w�ɶ���3�	6{ѷ����U��J�;�G�r�w������9�~�[�m
�E]7��
jK�)�8���s&����ߺՒ.t{2���1��A�R��|Mُ�I�������P��<p!~�xCB��K!�,[	�����a�:�e��\���o�������[3�auE"�FJLS�OJ�_>
�����B    IEND�B`�PK   �f�XK�h�� 6
 /   images/f2a2d8b8-8493-40f2-a2f8-368c45be6cc3.jpg��w<\_��;B��AD	�;A� z'��3�.�A�F�N�ލ.zo3z�Qc<��^�>������g����.k=.>n��*�(000 ����
 �����a�+O�=}����>>>!�sB""|���I��)((���)ɩI�)�10���z���).9!>!���=vH�ada�ab�<!��$�x��� `<���?���>l�g�x��O001�`a����'��E򔔙O�L��;9hR�3��
�)8��g�0\<J*jZ�W�98��ED����+(*)������[Y����;8zzy�����GDFE��MN������g����¢�Ҳ?u��M�-��}������ٹ��ť�-(l{gwo��q~qyu}���� `b�����!����?�'��9I��2�a��j�X����}F.��Wۃ�"����1�G�*�ņ�������_�o���� �����0I 2��߱��c��U8�w�ZH1�ӽ�.�"�1K�� ���o2M;�g�&�0(��]���9Dt��;�lC2>\��L0v��2x�3_pR(T�m���d?9��!��� ��T��lق�Ѓ�'���0I�\ ~YE����&w�v�Zr<�ᐪDC���%v��+�R�W�5u��`��W�O���˵ ���%]�r�E�M�Y*�b��v�IU�7��l&� �_���5����Lގs��q�<Qٵ��G�b}׵�Xɭ��z�ߧ��!��_����v?���((��v�5p���E���8�5�w߀�v����ᩣ�by"�/uD`%���h�)߬�g�滙����nL
J]3L1y6�ƾf�ɱv?^����~1)���o�>I40�������_2eclː�������ѐ�T�7�����#�`�?Z�\�[\3l_���h�ɇ��]��"W��9���z�Gޤ{,VN>��ɿJ�ı�U�;��Hs�ճ��к�n&���ܷ�~W˙�'
<�􏞹�
�W��$�z��~RQcG�r��gW��!A�=/��;�g�<�a���/"���ȉ�ա�������������G��V��&�v�85�m��7U6�
>��oiN�)6��^�?�۩�q\iP�Y%5a"�o��T_5�@��E}K���f�������!ӳV� �rbD�kw0�_h��]��\eKC���h�����j��c�7а���Y`�M�L���aw���F�A�<1��F]_ז;����Qf>�oP<�,$�n�o��%�S�3�ϧ`�n4�mW���DÑ17���VN[��q�����n��'"�" ��)�L�G@����C�>ǵE}Zv�᤯ͯ#��o��d�vEhNH�+`��׶���D�ֵI��:=V�~�q���k�W���Ж�d���c�0T�)���b!_�/r�팉��$Ex�X�)��ȉ��*�ǈ�1{�G X���jk3�\�F��ftp��L�K��3���|h��ݜC�S�f�{17H��(�ńI�"�y��'�v��H
�4��&��P7]�o�JD��u(1z܂W�X$<|��-����Z��}�+��s,?��0Yjp���Bt��7�h�,���7�O���_��y(1������ߏ|���iÆ=w�Gr5��K/����ڵ����34:��@N��U������D	>���oG6t۸��mW��B�����������~+�Ѵ�M�~�6��3���=�,�@�/�̫��yR�׉}�tn�vc����ټ�����3U�z��(`�U�#��ESh�X-�nJ����!�K8�L�I��ӵ۴�$�JJ�p�g�ud�L�������PE�I)k�~áPe_j�D���"[{O��A�[�&!�$�����uIMs�]���` ��D�mI�������-���ݹ�������T��
�X��&R�w�~_���Z`���%��A&N�f'.4�Re�Z��� ���\*Z��k�1�� �@Un�Xy�Z:���_��q*E�5Q���I00q��e����v:�1c�W�a��ջ����6�y4��7��f�9C�"$���)veZ��y�:,¾�N
��_�2���l���0�y� �W,�8����Y��=�����6�0&&��#��pp2�5 >	�[8�qk��X.����'� �W-*�o	!���Ϊ�6�7�Cȵ�a��(�y���&*�/���5��NN�X���9$�2��k�Q3�*e4W������C�tXIO���-��\K���'�]5�z�W�t=jW0?�\�҄#]�r��s�36y2*0�u��	�b�B�,����u�����f���aS��w;=_�V�����D�i�BR*� r\�OfG��ߟ�܉��"�8]��$t4�h�$r>�C��T��v6br�v�������l��N�:&kȮsy��{Z�|�����*"',%�C�[�����7�/V�E*=��rc�Y��,+�BW��dcICbԩ1Z�t��'��G��ej�~,&	u�bZ��r�%NO�/�`�����d˷v�A-k�-�a��
=��VG��{A�� �[p��I��G@���ڪ��0�R���6�2��/���Qw_���*�VH����r���}o�}��_赛����^�_FA��/�x}4A
�����`fea�0U�S�$9�����v�\�ȡ����e�K"/UW�*�\��H]����;���oU��Խ��#��/7��u�)i�\;�~�E���*�AL�_����D��[N���u�<�J�lזّ��I�M��U�ϽK��m��r��")�ޅt7K��s%�U�3CJZ/F�i�&�#�b��9xX�g���(yr�~r+���:����=���H?a����K�<�����g�t̓*����0��~MYW�v%W�� ���d���0Y8���	��E���|:��=͛��n�Yx�
T)��gG�	i�J$\�r�d��m���k��m^���/=�� �5��:�l��d����_��m8і��V|����9���<MA�VW�jso�jmר<���>���!D����!;��#L<��S�ڶY�����2���2���ケS���e��8��H�e�;��/q|kOP~wF����9����^�fvf�oة<笃����BC����S,�'�~�
A��o�.�TO�{By2���g��ՠ�IU#z����{�K�_��xnq�z��q�[j�Z��JM��r*�Vd=�6W��ӽ<؎�����!��m-�84N�����~tP���7���(��T�_�3\�@l����;-��P�~�S��qf��h)�o?��	�(�Np��g}�^�4�~V���r	-�o�0=p�s�v��ʑPf�U�� +)�ׁ8p�h��:o܊2-0�p����`Ŧ���@���\~\�Z�K�m�|=]�sZ�[�;<�p9��׋��,��Fy���nT�fG?79���啵C̔�x�L&�I����G�����iX�V�U�G�c�lsV���貪6��Nb!P<
��5ݐ���������{�Kl���@�:Fu�\�6)�x��_m�x�HQU4/����s}j�ڡkf/ekB�( I|����V��o����:KmR�١���|7�!0�5化
ϾLT��)5�[�1y�"`]m����C�?�_=Jnoe,ȥ�.�~�F ���	qn1]�O��.,��_��ov�����
�у"M�g� |�`ǕCD��;==#��9M�#S]b���a��ʹ��dR�+�����Α^xi���h
��'�6W{ �b�����g��9�{q��n7�Q�}�(��	���FK�^Ν2��AY�A�[�Xq[sz��2֚�Wb��������7}b{Z)Z;Jidi�&W/]'�Λ��to�zo�H�mL~lpe�qA>�8�y����uţ~n�ŕ��G_tĀH�a}�g��JŇ月�}�u�4�'�t�e���J\�'$�f%�`��;�Y�G@����x<�H��d����:��[����%������HHU��9������y��.�I,��������)>�Kj��%�;\a�T�;mY�N����_ՠ�%B��2(���b'��2c������ϥU�6�s����x�o���yH��b����e3������>��5�Á%�����2�h��E�׉��f�"��C�3��dd�(
�]}|���}\���E��2�$�P���U��r<(t�s�H˱�w�[��Ž��Mik�iPM8Ҏ[2�#�H0(�0՟qGd�Ж������`�RW�%5���~�r@����t�jhME5���'o��"�(Ͳ�/PO%�}Wr�>?7�"�1%������b�5ʒ�����+�
�VYa��܉��9DUVl�.V��l�T��g:����_	�8?����?"�y�3��6FW	Q=��~�y=�������W"U�fN���}%`=�D�����DN��vU���PI+�=�࡟�Jy-����w�BK>�x���/L�N��o��@n����_߬3њ�ZtuF1�h���K�d�).@���(�{ RH�i��{�D�N���SoP����P)�o�@��5!�!�A������h���@��V�5M^B�����q��Z�A �x�#�����r��8	�\�Ã����әR��vj�E)�@�v!kG[���ӟ������m����2_!l� ޳�6���V�V���q�!.s�4��%�������~#ɮ3d�{-U{m��yI���?晘�ܔ��PV���3��PNu> \��]��vB������ڥ.`�f���PZ4����ayȓ�p% ]Uʢ⫨����'��eB�Uk
�����QN��S�̞zW'.wF���L�_MϿ��r�*�*�s����'\i/�i˺��H���2"�S�ДM�@u� ��|�m��{��j�S���#���v�/�1S��ذ?��C�n<f��r�=����G�����*"U�e` �q�6is�#��Y�o�x��
���;�)侖�O�������y)|��O��G��*������[Ę�6+O��L�m%Q46l��l�T���,��H�]i��2�/оY�(J<\�^���"z6$��qه �����E*��t۰��[��O���C��L�7T�Td���+�?!� aǐ���X�X!�T� !�i��!�6�즷:4���h�ZiQŢr�S3�`����PqL�O��r������)yo�
ɘxcы-Ɠ����JtI�H�"�VܗK�pTj�d�z�y5N����^��J��kw��ʗ��@�h��U��|C�!2��B��ק�����;
�`-x�	N�߂"mQʖ�����C.:�S��2�'�]oc,�D����؈9�.-��Z�*&U��8@5�6���d�1��E��3�ж�/�RJg��;��;���%��&�O��*����q��u��_��i�V�����u!e�qڊb����-Nt�1­��߉P��񒲄�	�*�~�N:?X�d�!����٫$��$�,Ҡ����G���x.�6p���pU�C����ESY<Q��{8���Uy��`#��
O���]�Y'��X�'*��%�Ѝ�W>�[&
�*4sd�E�Q�K� ���2��� R��w3�\�Q�qje������G��/kzDN˓�.�~�����_��W@�R��k��1,�8�����'�Q84��IH�rS�6¦�D�F�P�V�\?d�hQ��D)>�� �lR�a��^/���^LS��8{Ԁu�(ϡ �}��%�o�<U�8R���':���>�`���8��<r�	�K��kP�����g�Q��ݘ��8ekn�ż�"&0�k�R������`w�rʀ+���/@�Z�������$�о(��Y�̵4
~;L����_���^��d�ۭ.��=/GO/pT�<SM�I��Ȼ�w��z�ک*F�F������@5���=�_5��9h[�n�g]'���d�_�5ce������e����Ulʡ4�U[�Ջ��G �ך�VS�и��
s،�� W����|gZ��A)��ԖZ����iSn�D^�!�g4E�Qߗ~��Oo��J���g���p�X�$���n�N"�6���O��C���l��<�䲱�b+��uho�`�B��JvkUS5�V)~D,k�����:V�p`T����h��J^��D�=d\�s>��봁D"^.��V'�?��xl6��@�w�aH�y!fFe�V:ZoJ�ޥ��"�d��qҀ� ���e�.�� L(#8Z�N>���+�x�������Nτ����>�v"Ⱥ�@��3����7O{s��Lo	SxOl(�,.d>�&��k����nex3�=���p��G	|NO���&c�g�����K���u�HN
KH�B��^�`}ʸ���p�0��z�L�4�S',�"�E:�uU�/bUc��X<շ���)b3�7v���A殾o�P�g��n�#���q�b��z�/�
W�����	�������zƽ�j��OP�0�a��+@���&����kO4?��D=8���$�59z����u=���O����O�lܞ]AT��:Lg�.�8+�m��f�����;`�Jk��+����{�}��N�iI�'�V�_"��j/en�-F�;��Tz�G�|�(M��ɓH��(�g���T��[tnj��"/��,o��o	@�����(#f��.F��AĈq-~����A
�N��o�q^����j��K2!U~�\nm�m�2\
*k͎��
���Nzøj}U"V�w�GC�UBǅ���yA�����p?2����4��l�^^r(bG�64P�u}`T�O���h�79z����]���=]����(Y{|�>�vC�<��0�5��y��^,�����ܗ�;��ѣ���1E�'ڶz\Q����,4>.`�LZ�a�h��Q��NA��T�]q�=W��
���8�mv	̙��r�q�u���|�	�$c��y��m`�Z�cj��r�[ؙ	�q�9$I�e��{`�O����S��Ě���M��T�As[�J$L6'�m�/ޛ�-4����PfhB2%
�ǋ}m�,���A3�_��9�����F���T	��"�d/9>R[��R�%��	�ȑ��^��D�fm�s*��o���p��[!Q� �����ۄW�|��˴�F_���q��b�ՌA{朝�w&L�,�ҩ�Q���ͨcl\��ߔZ�s�`���S[�I-�gh/vO8B��`ځ��@��z�/���{�S�p�i��Nkd����I�\�k6+`>ũ�&)~��9iƣ���`f���H�'7"���?�� ���9M���>�������%�i�:�:�����W�:�W�g�V�3r�"i'!�4T%��&�5g���>L�ح3���I���^5�w	72+����T�t��	��0�e��,&-�@��"�^�e�\"6�hR�;b�Z'�b󇲍	!j]������3�ݰw��(K�=�h�0�:J;�i��x6޺��ڃ4�Z�YBo�#�)����-:&���W���	�rh�c@[�/oO�Oy6d�:�_��QRD�� ��r�:�2$~�J��
��Ԝ3@p��N�v�_���4O�#V7��wW���;O�\��I|�Ӌ� �f�tö9!���̐PDm�����P��C�ra��N�qҵ��ҕ/H*g�����WS�\�	-�ťq0)(V��P��Y��?�U��E8���X�KB�XKٳ�I��ݜo4��������Xg?�.5�K�D�T���U�h�1ȣ^3�B��J��s���3��i��&�񋝺��ޫ ?���h�MMO�D�O��kt��[�$�5�Z��E��3f�f0�C�g�2�U"3���� *��nϰ�� �@��p��{HH���3��m÷�'v>���[�SD-����Z��c����@F�z����ϲM����Xl@4��9΢��w*���wo�S_���U$���`|G�j>#_�_{�������{��%���;3y	?�.@X�)�Q�b�?�@+����)x��I|3W|������8V�݀
��X�ͧ�
*�����)>�<8�бg���j���@���Pi�DP5��4y�+0�[�y�?�x�S��,�+0U�~�]�p7�����*K��;,����T�ęY��Z(��&�������$��񄈞��".�(ON'rHŧk����6��S��կ���A�ͽ9���m#ڵ�/���T���k9��8B��%��
-Vm?O�%���2S�ὃ�t'��~��Zj�
���&5��p�زY*�MkX1������U6� ���*)1�Bw�U{�o�H��x�L�W_�-��y�"&�a	�$�~��� *H��W�u?n��8��K ���r��D�%�سɖA��o�]���K)ŉ�3FyF���k;/M�0����[:���4�����Q���rg����-ū!:���2٩�(څ���Tg��_���@���=H�[|�j����+4G�+X��&�FL����9����S�쭙������̠��i����u�5���sǛH�`9k%��P�YP��MY[4~塕��+�JM"+��s�n*��B�o�W�8G�d�$wwWw`|�H�oM`K�B�=��
[\��~�{;����~6�ꎡ�[�#Y�T���\�\� �������ڨ���s�N`l>�j�.bnU�l46U�z;8=?O� X ��hx��7eq�F��l�iy�V-iB��X�lqd�}Lف��_�ye�L��n���rq�<�-�{�5�O��U)�V�՘��,sS��s�zњ=�Ϻ-��B��'��$���G�!Wbd�	�Hf�}ua-�d�_���}U�7�}Vo�{���Posr^������FL-t�Ľ1�T�im6�yӰ���%3��T5��3c\{']PmW����E_���0G$�Q�rdye���9~�
���|If���)�\�:$4�5�%㸧^!�a�w9\��K�ЈV���^ͺ�����j�n�r��v����C���&�8��;����~��$g�ޟJ֤��v�>�I�i-�o0Hh���dR��O�J�x��J�r�r/�%J�?���W��_���3G��w��Gm�,]|5ly�~0L��3./�2��X�<���2�����ո�`9�c�L�u�C�8a�vQ���E��z;Xm�G�,��\`O�߾c�]�ʵ:� Z޿�}��2�S��p��/��K����z�U9jAk^��>Ӄ57Y�����y$R�Hz�So<�������f��b�r��c����Jf}ڮ��\o=#�C���$:-h�UwkI���{q�"�k<�K&�=�Ѫ[A��_BX�"gV���ɷQJ�*�P��T�K�.�q����.z][t&�'��K_��-s���|�N;���a��ҙ���`�&/r7�.ï4���*E���|��`Q�N>��B�̾�E���5�x'5�[`�My�i��o����2�2�������K�G��-m<Q2��.�� ڕ٣�rf����Q(,�R¾�/D�>W4ж3r�G���0!��ܱ����r��K\���./�51�]R�s��/o�;�;Z�LʿjŜ{�`4�Bp��O>�����狃�\f:'����Ts[����}ԩ�F�R�'��]�������邾��l�*�uX� <zRj�1���}��BR*�ƽ�3��`��@G�S�p�mKW;Jd^�`��^3��ξf=5q���wGkAr�A�*� &�^I:r�sW���%c^?��J�V�Mi/�e�:��@
T��6BeKr������'*����t��,�Vǆ}H���z����$�;�H���	�&�'���5f���v�T�%����;�i_3b��b�a4G�l͊�jBqn����%�&�X�~��V�<�S.�4�S���r�k,��v�GlEy���G�TI�B��+يR�j�U~�3�Oiqo'ZkϚ�Z���x�ѽ�i��w�щo�/��^��w=��V`���@�U#'����:1�:�^q��P����k�2C�
�D+QʒӝL<�Yg
;EY�E�W��ùә,M�#j�Wz��isp0���C���1���٫W螺���ݫ�2��DE?�e���,]�o�MՏV��_�E�W���K��8ծ�j̺uK�H���j�L�f�K5:H�O��r��?7M���^^>�0�TO�iUg;cO��\
	�l�'���Tn\�f�2�U(��ô�۴�g������V8�_�9a�L1dJL��jq�Q-ɰ�Hfk���6!�\Z���T�8Ǚ�\Ld~���xG�;��4Y��ՈMŲ���꿓�G���^q�熯�+��Y�	Yq��h�P�
_�e��2��T�:�o_��/X2f^�)�w�߽�q��|�L�OC���Rt����p���e�������9��W��+�C	��u&���D����q��8e��b��d����-2�ޝ�-��:Ľ��[���#��B�z|�a��퐗vTv'�F4�&y���wz�\	/@7�������Mf{.P���0�#E��r�@�&P^9Q��j�^s�B��OE.�����#�C��\@�B���x�+74s��Rn�x��n���a���v��J�GqRc��� ����x��0� ���V�G�)[��tg�%���9�x�e��-L<��4�Dkkmlʷg��p�<d�tz��w%��kV¨�>B��
�IUM�d�A�aq�7��3�
m�S�/�D�*.�o���Ű������x�L���`2ԧ�G@$U�r��JP*��	s�0�a��7)���� ��1Rm�/��˝Y��韀�# �������V׿��l!-�K��e/���"(	*��U�"wDѶ&}� ��F���Y��ӯ6�ϥ?=鼭r9Y���x���6Ѱ�7�ː/�އ�j��K���S���Z%�6�J�vDHVZCY��w��Y�,����+�����-sZٶ#?q���~Ň&rmG�܁��m������������6,x�}�ُ_���o8�ug�쏋���[�j�wY�x���g��B�e��Hͷ��y��_��jm�Dª	�=.��E�(#�W�9r%���z2X��n�$�#��У�c���ioK�^|�����o(��t�7�@����~�1M�<HDw�f�Ɵ�no���� E���<i��g��j�x�O��e�ScI1���d��@�(�ļ����!�K�����ZF�m�ģig,��\^(7�Q��������3z]T�<DV2v%��0���Y�+<��6�eڮ>�(�v(���2��0��CW���9]{��D�w�O�ԚA�S�(DL�-f����wo��56ٗҖ���P��*0��/����,�PA������F���$5ߩ��N��W��(�N>�ʀ�ǧǢ�Zt���z&u♊����_�H��s
�O]��f���G	�
H��&y�GEWA���fo�\n&�}?�BdsZ���	����hv��u3�Իmj�-�i�����1��������'��Qh6#=Rvmȩ�Aw(L�St�mMk�^0�����[�X��䝙��]�Ԥ[�� �\tC ��C? �W�H#�U���(�T����l���&ȭ����_Vl�N8*_�c�Ѽ��7��cqI�&�;őy_�j��:o��J��Z̩������ثD��񌀿X�7�5��v%����K}�����a���43�]J�uA�,:�ݕ��{8�|`�t�4*�n�I�<����ﳡsQsC�ꑷ~�W��Y��v��lC�Rc%�q�p/mE����%ԕG(�@MY��6�>��Ӝ� C'�B�U����߳�$[Z� ;l������^ۃ��s��1�OY^�	����'�rf��D2r-�6��
�Oh~�*1���&gH���:�hA-���4�����4�#-j�~��g�� �L�\7��/~\�(��Բ��� 4p�+C^���䜞���|q�JV>���:o�����/1j�'���������u�p;Q��VAYs$V�<m��x�9M�f�b�n�,��߆U��|348ϟ�#.G�l�i\��Be�~x�N��O6sLH��UO�x��V+�`O�͈=O���J�= �<RD�뿉�xʇy��$���J�Fxv|�U��z�hu�.}Xy;(n -IX��Lu��B��.���fۮ`��CTW�������A���m�ML��.z����*����_��#U�0�ӷ��_,����tI�o��Sr�,�mS;
-Jt\�3=��w|xQX���&�ɒ����v&f�i�������2�Mo ��7���,����~pW;�חCO�9�	cǈ�0���{^��f��(<�i�ƺ�[�� 
�%p�ek��:���h��-t '��QҌHM3&�K�5%C��q_~�/?v�Ď���K�B�dR�<Fx�#{��E�<�����"D)j1�Ҷ�H��k y(�4׵��������oeJ�8<ݍr���p��w�O� �i*Dq�'����)H<#��UUX-���ϓ�'
Jg���&.��Z��gͰn�cw�,-�,�ߴc���k��^m��>3���'����v��d������f����w���CX�����3$v�n��'�o��z��b�e�U��f����weQ���G�a�c����6�%�x�c�[{O�����I2�ħ�0�o�*sl�w[2ꟙ�p��� ˖H��0)W����^��]z0:k_���M��%�#m�yh��-h��[ݻ�t�S�u�G���)v;�����60�Bϩ�O�zKl��Hc5:�["�z���j�Nb3��v�܁����Ԃ�?�1��U���]���Mz;�m�g(.ׯ,^�i�������2�b6/����+����e����<=�r&�!�_bO�zP�e�޵B��&i�P�Y˽��(��y03b���
+�4A��G��}��d����E΍�)B,�M7\�|�a�=��%R���Hp�(��[M�gC����ИL v��]��g�%N���3����>�W�!����"D/�9w���z��w̓�Tx��"�/?�d�r��+dx�Bf��7��.��
֭����Jj�o[#g��f�m5�dq�ʙ>�ְ}�90�"r��ǁ���	�/s���1�U^)��&е�Z����y�i�4�7)���#���s5޳v����	f�-%~�dgwnC&Z�:yRR�o%��A<ڍ_����g��$�`��d�k�L?`U�7]��܄΃Y�w�Q�A! �T�,t�9?���5 �Zr��70�t����tQ�qr̡�֪���Dc8�2sX�s�L�zE��<�<���*�g��wJ=cÜc�_�ṅ �=�/b�	0���E���d�״mz�ι�m��Z�Yg�t:�{yC�WR梟���d�?�ఉ0���B�!6���G�G ��-��a��}�D����sO��&I�`�F�5\�*���$.�o�����317�9�"Y�|��
}+=@�2�/�7o� ggd������*�|�dC��艆D,���|��������E��r_�u*Dg�V�j-ES0+�ц'Xda�'���'Q!��F��'�IydGR�k�kl	��j���e��������U�����zqQ�Y���ǚL�^��uPL�!Ս˸;벾��Q�ݽ"1�JbB�p@z�����J��[��R�U�=<�?{͑��)�7]Q���
Z(W`�ԙ�PĵiG��z3�[K��Ng+w�Df*�.��h��z���Z9� ���L\\�Ϟ�e�K�5��@^�,���-�J(Z7�׬bp6<4@ѹi�\��,QT3T`�q]����AF]��>�u:~0�fo�o`憯$��w��=K�#�ƼtkMN�e�5��b���h͈?�9#����UAN�3׊��dy;��@�a�cI�H^��H����.��9�S]�H�dP6��Q)-�����@��W����Y$��3�ڴ�-�OȪN�((sW����䂰�CC@ǳ�1��K�+����7���F��h���o~�������N|p�]TQ��c�P��Ǳgۀ�w�� ��u�T�2@�ˎ
|L�����M��@�H?N���`�Z6���6�g9E��5��=���Kώ:���������ꪎ�c��n��?w�#��iP��c�J�޻���:��sJ韞6�[�Wa>y�T>���S� ��A8 ���{��v'k�Х��J�|��y��tw�"]&�ɹ�FN��L�[Ϙ�Or}�T{q{v-?d�e��U6&?H~-̯3��cs��z�#9?�;bHB�j�je��%ɂ�ލ�oU��2_���C���e�	�c�U��53��'!~'j�Ee8MR�l�g0���M�02��`���esM+�Rh'����z&�aBK��}�G�D.(E����+�`�uK:��a�����d��(��g�mf��	_�GG��2H��>��=PH�B�����������<����ъ1>�V���,��&tB���z�P{2�:<ȷkV�c,&�u7} ��[�uf�l1�F���J	M)E�:�C#�i�l��C���b�IJL݃�{�h�E��L�s�5�T��^lR莌(��I�tC��*_�2�+�ǣ���̼%di����T�տ~P���ؽJwti�.^�4'���P���[�S�������ۛ�AϹ��}��r�ˉѨ�.�;�I}/��9��%�Z�Kh�.f$������F�@=�^`*���J�I�daA�3s���n���M�j���o;�3�+0���k5W���F�nǷEJ*�u�0���{���s�wt1�2��!�s6 4�U^��?2r(�{^d0��V2ɕ�d�ɻ僦��)��묏�0??5���#e�ɥ�~U�������C�{���͵��z��؀d:���ddL�"�ْ?�VWd}]5�(�-��p���
��n,������-É�@� �{�PO�ڟ7JۃqM5�l _�O��䩖��~�(�N�.t�`l�-��²��(z��W>+�z���P�z��#��ۻZ2�5�J�?5��X�7��>z/4�u�y��u^��)"�>�E}X�pQ�l��o�0�?c^�)~���N(.�mΞ_�~P�w��F�f�U��6��s;���������78���,��CL�[�w��W_����Z%�ERJ�A���`K���Â��&(�����/�3\�;���}�*7���h-��T,��������ѩj���l��k��Z�x��f"ph�O�F|pj���E��|��D��yMԝ,&i�����,_�m�?EF|l�[
,y�:��{�X�$;�壯�}V��j�ę,�GF�^fIqCj��^�Y|�z��M� ��G���9�|Z�>4��`y�d�u�O�'���~�;�ij�j_��E֝��8�:��F�����/S�t��|o8�����#e9u��x=~\Mhl��Ī�i2���{Y��bt�-ZU����S�����2�diBι��V�4ˎ�.�"�`�2y�>׶i��{uo�HO}f�^n�"����X&���1����ͦ撕괷����g-r�9W���sz�<XЮ�D:��u�:qܛt��^+h�VX�ai���U�Ţ~��b��u��n�}B���FCf�$�1F|g���J/�7����@1xo/>.Z����}�W��?�s6]�X��c�%��F�ɏ|P�#7��ti��M:��s��/�tdęŁ��6�t��{>B����Y�V�ňه��q8'����L��`�"�Edj��D��iH>����-]��{|�H_@�B�������Io;����2e�N7���E�	�Xs��a��0��d��&�C���>6�D��%�;+ε�L=.8.�3�*��N?�|�-��+�\��,.B��#D¼hG�|��\�9[�/p�$v����9ռ�ڗ��k�7�ޔ�9����gå{�SS1�z��%8��`�14Rp�E���7r_/Ԛ�R�i<��h�`ܔ$9�2���C͌���}	�v�&���a�a�O�m�]B��I�U�j��z�?r����"�(nC��&$2D�8�4gX�%�^�ɜ2�2Y͹���v(��d�2W�������_ P@���5��uo���3��jB4EV�v����߿�~kǥ��we;���^�6��9�\�v� x�}*B���_�� g���*���� ʳY,/f&�G(;eFYAWRs���]� >�xoR�g�����T�]J��1<%s�����G��~K%����c-���cnI?/����� ����{j�F�?O�+��O��|5�Y� h���&o&�;�x"idQH��1�UP���<dׄ~�Z���>'x�W��(�[/���qnwƫ�2� c#���t5�w,@�or:N��#�F�Ǻ���yR��=��Z��<�|�/揺?e/��o�0���mWBo��	<�X�� J���z���i���\�7n8�}���O�?������~�>Q�On��rrP��u�k�
x�F����u��Asep@�g���䫩#k�=1���J�S�U���g�e8�y�4f��{�2	>�{��u�?J�[jZ"�2���JpC�#��� �[��L�		c��$��U����*o�J����W+E���A��M,���I�+ͅ�j���n��|��z. ��j���u���]�)�%P}=��>)�S��i~LSy����;t;��I�� ֯��sigaG�����Uvi��<��>!����\��%zP�������� �ۛ�<ۛ�V�i$�$!� ?J����ֿW��t�Ћ���ºįj��QE�7��ҝM=?
 �O�~�ҾP��.~ ,��C� �}}_/O�� *�7��b�H�?��+� �9�>����Ŀ
uGa���|L=��z~��OxWPT�wZD��  �5ǡ?�x���f�\�x�e*��:4�y�:p�CV9
��Z�
�v�Rk��<�w�����h� ZƬ5�����o.�� `:�U�x����Xd��$��n��#��T�����x=5<� �,�|���j��a�pT� ~�W��x�Ht+Amk#!�ؗ=y�Rzu��d�x����bx�8ڑj�ŏ=��5	��sp�b�^���q����P�-�᳥[ʷ+3�;I� Ku�I�n��ua����Ҹ�7�����O�ax_K_�j�����?��5�!�3�<׶�y`���9T����>�O_im�������:�p3P%׌��UfQ�45��jϨ���a#cDڈ@��Tc�GW��#\��<�����)�G[��u�8��]����:�U�� �G)yn��w��� |��O��G+�b	*	�n;�'����g�K+ˢ����=8S]p�	|Q2����t����#H�^��m��J�c'�WN���>�fG�:�~+ʵ����P�f�L�엑F;�]�:��J��Rٝ�9�ۊ�Q��%*ַ(�	�atn���.j��m�q�	��H���[��ȟ~X�a�NH&�oj��h�� �\��]��&;�V��8��f%
���?Z�F��	�U$�e��x���6��i������;�^������/p�p��I��� �q�My����8<Q4�#S�6򱴞����z�eM�a�5���f�Tc��g�$����G�/!�ϸf݁	���:��>&|B�e���5������Q�[�Z��`�p~J1��ϟ���_�4�R��(GB8�S�S���~)�4��5i��Tu�-���#�֔�~E�;�U�nx��o��>%���񦻩Gs�[L���"��i�r �`�6y⼣��όڷğ��G��#Mm/��A p66x8 ����^"�&K-?S��	x���b�wt��]O�|I⫏	����70+fTI$'�1瑜�҉bc{����I�M.Ii��>$��J���weɒ��F%8*Y��A�^��� ��,�~0xKF�\�д�RݢO���
���#���|
�}��^YGhU�=�<��� ���A�֧ǉ5� 
|]�m���]Kz�,��;��L���랄��S��e�(��T��[���'�χ_N���}B��1v��y3�Np3��1�wj�>=�9ռ���X�<}�L�Gmi%ڈv��G��>�<u�����YaMD�ѵ)>kXu)<��@F�n�����?�CQ�վY�i/�r�V�K���l��^�ܥѣ����>d��>$�Yi֏��������0/2}�;778䞋��o���F��,<G��5��g�0sR���8=;�Ҵ|'u�~ ֵ�=���Mϛp�sj̎r��9Q�zt��k�R� i��6^�N��$��ȒIRAq�ς�>���������;O�?�<O����ƞ&��Y���`�[���˸��H��YS��WM�f���^:���0�$k�!B��ѹTc�'����:,��)��Jo��X����_�L��q�V��-h?��X��U%��l��l��� fm�wg޲����_wF{O��cR�h��3q⛭eb�̒��rJ��x���{ds־c���"�O���c���+������1�]���v���Eg8��о�)0�.�_V����W��R�L�01DKjg(���'�\8���������O>_��wӔ7@>��:T��Z�J�r.�����8�U|Y��r�im�&�ԓy*X��h��~��o����Y'��QDIĶ�#i%J�|�$�\q�	+�����j���h^4j�j����۞nqU���֏a�,�����\ż�K��bF��I��8��U�xt<�c�j�C���e�� Cl��A��*��y��6Y^���/%W�84։s�b�����U���|H�
��� O�W��E�S��0O��o�Y�^�}*�����^�'Lq�{��|J�Q�X8���� 
ɸ����$r��Ep����?�T��u��p���8=zz��MRW���V>�����u?��V�lw7���L?4�Y��P1�I5�g��%�|?֦�<O��h:�`3�_Bbp��>����uiu/|�Dk4�kv�� ���W��S���Chm$��� aB��'��c�[��^�h��P��o�/�>�F��_kzޛ���6��ܧt?�_o�������'ß&�v��ٹ��6q�2?:���W�Y���t3������^̩�^A�
���	��	'�����c/�>���Lx��>0�ͯ�,<?a<v7�i�JDȦUٴF� ��6>��o����V�7�5�H7��Z0�3�,=��k�U�"���$u��}~���|W�Bx#�����]�ђ{[E�$,1��]�,`0!�9 ��1���8�8�1T\�T�ӓ����)�'e���'I���BZO&��G�]�"���ӯO��O���Q2`-���׵K�y72٬���1���>�����\xDh㳰�R_���~�m��R`���vK��� ��!�q�W�ێ0z�{� �w���6�%��F�<X�-���LT+��\������
m\�n��H ��^��ܐ�T����oj7V��i��p���i�3T�2����s�b�o�feO$q����K�NwU�9&Ty$r�Q���\cJ�����H�W�/&ҧ`[��f�Yy�޼��9��x��^0���|W���k��^e�Ɔl���'�ˌ��{���:����G���;S�ba�k$*3��8$�������\�*�y_+}��zs�c�(�Ka���ۄ�8��?<|�쎜��4�y��!�9r,�,�һG;��o��o
�F�쌍߭1�����̒=�._z�jʤ�#�R���j�!�櫣�VR���LBy��� �N�����?�<���(`�d#���o�� n�e��_R�m�YP�P�kd�i����X���j�ƫ�� �M�ψ>�o�[��:��I2�3�� ��t�K�[�&x,�ʩ;y9���� ��I���=N;Ww�������������K-�̤� ��P�&�h?*���[xq�=ɞX�ʉv�0>a�{烃N��|��@n�4Ƹ���}@?�^�7���"�5�#�JC��^kY�9�O�դ��/�g��Ȇ!��*"���Lv<�.U��p�x�x�9��V�7,?��T��Ö����ooR	�Ӧy���~�nǰ�Vuχ��5�]V��La��wx�u�23@#�n'F��b� (��~O<� �*/����|��H��X��|>i��X���F?~�d�Y��ȥ_�>hgF��9Ɍ�qK�@�۔��o\�{�(�F�1�Ӷ?���2��?:�H��i�)-[Px V%��#(�B�5:|1���X���D���pGjd�͖H�6��g���D�$��Z=� $���C�� �� M��D����%��p�%��p�@���מ��t
�fmc�E�5;-kDҼ3��鉨x��H��@� "�q����{�ɨ���s�ZH�]�|���^����@d��n$�c>�����<y��Zǉ�o<�x6t��I/���m��d{�h��ۺ����f]?�݌S���������7�	qt�W͔N��������槙=J�g��|�>`��)?����f@F�������'J��i�[h:��	�	�2����#9� x�+V*FC�H��D
������TWWlX�[�9�!l���Q;X�}�@��â����>8�YF��?�#JB�e8���J��df'9=�JW��'�q�=j�!Hl9��49u���V찣HG͟�t��4�4�t�6���X]�Ɛɹ� ڨ	E�Ƕ=*5��;�G��e����*M�Ѫ��+�\�y��^�R���3���1����G��M*�˴���G+q;.9 չc�ݷk
�F)��g�WUQ�%���4���j������ d�Kߎ3�Jт���94��^~��«/������1�Dڲ|�=�T�7ў2Ú��7ß|X� �<�I���[M�D�E�Ig!G_Z��>����ԛFõԎ�N�zG�?e��>�/|Wቼ=���6��X�P�8#7<S�� �����񍭥�
̺��������j�����yLq����G�q�׼xe�ot=6]>$��p�\퉲A ���k��>x���V�/�.t�����7���vɴ����OZ�}#��߂4�ĺ=ލ�[�%��\J�$�������Z��[�����9�ކ������/�nF	S�Sة�j� ��|}��p����e�h�#J��^���O�A�Eo��!�;�A�'��kx~�m.$�2<o0�a_w�ld~�I9AB�����c*ᤥNV=g�� �%բ����&�a3Y����K�������d�Y4cx�k**��r�x�|a���+(<E:�+j�{���\��F�=����-����et�}��5��2���5>�qf.�q�=GP��<_���4�hr[��)t_6P��݀�>��j���c����מ!��֮&hؑ�1�Ǧj�����Z1���2ۓ�f�Q��\��.�K3 _��Gp+���p�;*0>�V�#%Y��;�4o3�d��}�L�uk������� b�� «�?{��G��_B�޾�2n)���04�$�������#t�)�H�(؉���U�'�-��p��=������{�k�ڝ�����?ֱ��6|�y�u�j�}�Q�Bs���:����9t�!��^ߝg_ʿl�0?�X������ $�q��I$�����_x�_^&���\A,�c�#����ں�c^��í&4�K�eh��|4��G z(�{�;��Q�
�o�r̠u¯�+�����*s�\��˷�����Z����;�NU��h>g��%����Y��`�G]�Ͽ5�M�$�ʆ'�V0�tzz� �b�_E��8"�(׀�����?6Gs��{�=I:��D�8*�썄�-����#9����7�!���܋��F�j�.J�:ӭt�]z7���kKY�!�D�b88b22:wSMI«��f�� ]|Z�ZZ�5��`�wt�H���9���1���]�%ť���7���H���Mg\������F����	*��,�$3BI��H�a��;Z�s�_�1ئ���_��V}�veD�<A(W��N3|���*�ҭ�\�WGؗ��Q�{A��ڍ� �U/�R��Io���c� B��!���|G�9_�nт)n�K�����(��]�؁8����}���:3�y}����|�r��,�����+ğ~x>�MG[�����Uvf�TRY�_�� ��_���_�:��&K��@ �?1 �O5oO�L�΋u�jQ���12C
#jR��rD �ɢu)�^�9�t{��|u�� ���mB"�V�V�Z�&�*�27���Kot&�ɦ[�-�%���.HN���_=��_�<�?��l�>���j�w���U;O��+��ȼq�I$�ֵ;�NI�3�������}+�SյoR��E-�}/�|B�q������o'N<���X�a�@��r�_Ư\|Tҝ^�_
�Ȑ]��+*�d��'�=J��/��a��_��Z��� jren"(]��{�5�������L=.Gx��}M����_�+�ش�Z[�'٥7��2�s��8��P�-!��G*��n����{����Z�����"���4�F
6�צ?
��.��X�ps��yx�^1�?�$�]�m���{Yo-��V�P�^q7�x�+�� j[��=�/�5	4ۍq��[��B�,���VO�!�#8>���M �9�|.r~\�y�E��Aj�/�,�d2�\�M<$�N�����t��J������'�<O���?��٭V�^i�d�Kl���.fl����/�^2���ѵ�Z��i��nd�d��;_d����c����m�nF�[ϭ������푬��E�ӿ���k��5��g�O�+׮:b��"�W�>����[�����˽B��[?�QB	��N�d�3�Ȳ7<��1R�z������c��ƍ��b��� 3�[:������jWW���g��T^՟����y,�t��[��'��W��y�>vY�n{E�[�{�Ax�����O�vQ$��<��3��tQ�� ��Ժ-��t�^�>x�YO�٤��eH�fm�J��/8�zo�� kM�>�� �l/a�"����@8=k�����<,�|-����7�'<�W�OM��z��s�N)ʯ��?g�x��O�D|M��#P�ў�#��H�P81�'���*�M�G�f�'��`p�w��ƽm�n�+��Ӕ��$�N��|��;�|a�j�^�V�k�+��bl��8�"�9��Fe��V�aNWw6�g?��ig���ɸ�;U�8H���v���-��M�-��o�t��bvn�i1�A����D�Əi��B�.4=^Gf{X.Q�̤4[�ç^A��ľ���.��xm�?a�C�yD�0�I��o^G ���ש��L(K��Ϣ~2�Q>�B�I��ue$b�	6��m�g�g�Ď��(�$�)ʹ����#��Z�m����D��>�ykm�-ĳ9�P 9�V�l�~��s�۲Y�ły�� s���^�z,��Æ�Zr�Fv����$,�*u��QI�w�쓓׎�=�Mu|��'���WD?(>���
r�<n����q�L�֗�'o��µ��MM��Ci���w?ʩ\���~�ˌs��Me#I �U�n�/�ÚH��۷�S�H�)��}R�u.����V��G����|Mo��(�!����V� �Co+*Ƞ}�-O�Ȥ����ea�r�`Un��{��I� 1�O�k�I����'Y|"�����h�r�:��ŭ��o�"�޹��۞��s�7� ����5H��k�GQ���-�����y�e׏��� ]yg��ee�o���ť�ŗ��W���&����� ��=��� ��� Uմx>�9�l`Ӣ�m}�Z�w1Uvp���$��]�N1�w>�7J
/V��=� �!�xY�%���BK~זZ3��$*�)Æ#pf�'��<Rxg�
#�7�w�=?�>
�+�xt=����[\G��`�,�l0>�G5�c�FxF���S������3\���q?7��ˏN8����4����/x'S�i7�p�Q7d$�T���vf��'���?�� ��)�~�+���C0����XD���Lʇ,�'�W�6>*��� I��0Sӌ�دӝw��?io�+�޳e�_���N�r�m�b�u�Ȏ"���ǡ�e)���<r�#�P$�w��v�͈�q�p��=Cx��<D ����`�>�׳�� �z�Z����G�΃}�-#P���7��Ί�wHXr:��/�[�v���si^���i:����͠�][�bU��n���˗R�ϙ����Ku�}G�o�r����� �'�\� �x�5/��.��߉t��7Z�`��m%IP�AAJ�T��_�?�����Y$6��������iV0��4J��%[c�9�2<'�2|M��5۽_C��}6�F�>I5i
ʉ��5e�6v�������ӛ@p���|;�������������-�n�ՎNz��q� �3�3i�q_��xRg�a4{�%d� �u�nz�W1�O�ƿ�g�y�R_�i������z��#�+��!U��F9��>-ǫ���A���λ��ŵ強�r��08 �NK��h��U�&y��b��?4ht�=�~���MՄ�08l��EӦz�y�����a��|3u;8�+y2��X�,u��ڽRo���� ��!�������k�I��Y��M�/nA�癴du�9���(��e���{�gZ�,�<F�Os�H���xq����(����v/�&�ƉD�m��z�C��#�ϧn���p��>!�Ͽ��&��ivӪ]Ŧ��5��mW*�>R}����;�=S�-�x��z�������m&���YNV��vpp ,�>n�����$Կ���׷��f�Hӷ�\7�6g�8?x����S�@�yv?* �]����9���8�#���2_�yO��X�\rs�\��[�+n||� ��#��)'�$*��Y\��)*q�1�'�&�ѭIG엃�%���r��YԬ�Zڧ�.Äm���g$�� ��/��������'N�f� �n��O�LO�d-��s��灚�m� c/xo������ݔ�1]J�g��	
�Q�yT(L�����גx��?Ѽ����J���$6R�u�hؗ��.Kw���5�S��Л�������g�����[l�E���o4�<� ��0N����k�ω~=�5��
Y�Y�P��c �$.3�J�°|/�|f�ִ�����Vр�K�rg�JpY��ڹ�t�O�1�6���%��J�n�
@'�޴�kndέ|I`�JC$���ȃ�����뚩.�m"I
[3��
�"e���X}ěI��V@�Oa��V$��7����>WQ��ζ�&�iHѤ�U(=;b�������U����9�[C+���B�m#�:e�2�nc��d��?Oj,��� ��mVIa�.��� '<g ��Y*��O5#���`�0~���MZ��c�����z�<2FR8��O��OҀ:�u�I���P0E����֥��e��� �� ��!p3�A޸�;w�s��&}ȥ�� ���Gl0�>�m=}��Y� iZWŽQ��������i��V.���_�}������u?��g��{خPh�Э�;���l�-�q_kvGR�$6v��{u4�P�.�H (�S]�?�ߏ>h�����iQO��=�6�ͧM�O���l1ߞ9�E_V�>������W~ӾYy�<[�X^�X�qHHIZFg�@�8�-�>����7:�����Yeu�Y[I���PZIȑ<�y��@]�ڼ�_�/�x���?���c�2A�����ܜeVt��0�� mʎ���?��>=�ׅ�5	t��Z��4��˨M�ώV=���o����NȽϔ�[�.]-���6�YٌF���A��v�k� �Ae�s����4ω�O�x�[З�G*�u	�yaeZ=�T���5�x�?eP1�wӯ��᪹,���� �N_��>����é�{J��-c��;ۉL���o	��隻o� ������\x��v�I�����DY�}-�V�~�	�K���oy���b��*����I����ڶ��x�K���'�}��O#<�� ��_A�e���x��գv�W��	��,H�<[���M�ˑ��%� �a�J�A���#9�\��yB�ؤ��ٖ�l�v>����������?ξ��uU�S���_�pV��L��7
�Q��Pv��3c��U�� ���8��~�W���e��b�E���7�g'�WԮ.l�k��yvlIJ����� S�n����ݹNN��	��BO�G�^>w�$F�m��7y|t��� ��_\9m{�JT��_�7]��uw�i�q��,~F��0q�ye�*���[����?���z�������쯋8�<(p3� �� ����� |M�[�g�������4�ss<7r4���8�5�&{��t?��M���������KiWl�����d6x����:U���S�����{�3�����9=q��
���㍭�ׁ|�k�vR,W1�G���C�@� ��^��k$R|0�n>�n.STI�S�����\Wп�+_�8|�㙾Zj���}�(Ǜ4҂s��v��9�G3˞__�7v}���)���~)��˿I��Y� ���ɵ&�"M��4�����F��0s�犼}��<?�mSS�Èϫ�q����̥�������~��>��A�x����,�%h�h7�d՛KH/g� T���HpUz�NFNI�ҾxsO����c�7��x���4��Q�bH�e n�s���\y6:�WC����~;M��R?�����!:����e##	��'�5�!��>�V���>�t�z�o�L/�"!�8'�8���?h�?��e���C{o��J�M�^�SvYY�/]�~n0~���/����g��?g�;u���l�
�R�e�B�I�I�j=���68������܍cA��A��Ko1��!%�	��0�c�q��m�Wk��e�t�������Ϩ�*⭛���Фq��پ\�X�䏦)�26��æ��1��a�rǑ�-�f�߈4�70_\4�ݾ8@el��;��OZ��h�u�:���SC%����gh���~+�� f���f�����і�����8����j�G���[���	x?Q�H������<�j���l,q�	��ko�!���>�j�>5��o0����M}�4�#��@�-�����s������k{V{�7E��� S�ߜ��T�v|T�a����.������[�d
O�;����3���W�v+�� Z���]j����mڊ����)n�#�%�x}�Y2�V�p}=������U��#��[ɹ�sq��W��� ��˵� ��=	��� �%o�I���	GVK]ߞ:V���0�t,��6�s�2*eOMͿ՘E6�o~×��|#��%eA�L�0�dg��љ�:q_/i�ǉ�tp�H�K3<��lh�=����|b�5��+��5kvn���s�wƳ�J��`�J��>�FS�r�-�k}f�q5��N�.��8�:ꓥvE�+����)�H�)OJF�L���w�?����G��-O�0�� :�=� ��U��Tq�%3� >�� Z��6|�}�����BՑ�� �Z��g�?�� ^�uflo��e����"w���� 1^����:�A~`�R��{0�s�|Yu�3]GÞ4��9�r�m�*�rFвg<w����GT���͕f�[qi�wM�B�lMі�7b���NI�'73w����MIg1��3�q�S�� ��wg<S ��g�?��Vr����W2#�$O�������1# ��Nk�?^���DQ��JǨ��H�1�ֿ9�O'�F�����݅~��)���a�fר��W��	��Pvm�p�S��ȸ𮁨GR�6R<C1;E�#)��u�'�����i{_�v��� ��<_s��+�0F3����{�����������⫸��aŰ#a��s��^�W�m�5��/��k��o��LĐN��z�5���'�[#�1m5F�?���e�]x��2M%˹�(���� �[�N�zW�wZN�����Fo��Fw>�������b��6��U�m���?���I<�W��^N'<eW;�-=Z8R�$��s*��6�Е屷���q�to�.��ر9�I�+���͢!X���UitO���\�sY��6q��HƋ�:_�C���v������u��m"Ҭof��($Kip�`uB1�����ae����5Ӥ6��?e����'�R����羽�kB�w]���y�����J�Ibs�=rk���a��l��+��F�umyI6�� �k�l7�BA��J�z8�kc�k4��J�����X�԰:ʱb>��\�.2i�������i�������X���#iFh�q�^3��G4���q��>%qs[[�L��yR,�e˰8@�:9��^\����zb��ls�^�'֮6����ɶ�r0��)�~Ӹ�S�����#u!����S�a=�pOaD�Z	�K&:i������q�5�����A?u����T�Q����T\�v*�ď�_��L{&<A��X\Yx�B��-��,�����dc5OI�g���4��mn�O����S����;�B��t��v��@�Mg�tL���q�sZƤ��-Q���i��q�{"���5��UL���N	�d��V�RY,o�'6�nYs�>b� ��q]ǀ|m��W����mJkc����72s��՟�� ��_|?�_�v�"�/uK�EΞ�;��Wc�)���G
�J8����i�t�1�-cc��Yn����$�3cijӢ�;�r ǯ��qY�����2�Yݮ����{;�V�3+c��:c�Zڲ�I���r��[����댡=bŅ���+�+��*Y��u����%ǩ�Tmi0� ׭+����Gl՝࡭�v���8�G�D�ZM��H&&c��<��ڥ�|�	9 p���F�X�l_ޢ���d�h����~����:�O-[R�R���E,&Bp��#��s[>� �g�2�&���C��6V�_ES��Upk�=7������� �SI�e���E��AR��8��4�ۏ�����O��E�<����P��(Tw�f�ڝ_ŏ��F�1�ڶ��^��bi*���X�?B,tY��YЁ�Čc�?_ҺmO�߉<mk*k�W���I6ǯ�`����.0#`;����>�F�fRP�(�C�W�/��B���f���>?�_���~���g'����_�߳5����{��t���{b?ҿ<�����Tr8�+V��6?C��-��{�z.�����<1��c0%E�.��Wʿ�Q�o��!֦�Դ�FU���E�"7(���ݰ�Ʈ��:��Q2�[Ke�,Xy����⽋����$��a�"l(8���*�����C�v���=3�7���S�|B�����7~`�YH
%Wڥ��p�z�_�~7��n���^hwo��h.�(�s��#�ӟZ�ۋX�� ��0�o�;s��z�	R�1�Ű/����Ny#ֲQԭO|� ��|Z׼��g�Ɗ �׭.WT��X�e���8#r�͑���~��� �1G�j��d�mŭơ%���i1B��S�L��sߥy���3Q��<e�;|%�Ɨ�K@[�;�c�&p�����^�~˱��W���ߎt� �h����i�.�fE�*��3����*�o{ak����3㏈t��:;�_k��WSMgIկ-���"�Cqyk�����\G��o~ў&�qe�G�����WkH�H���@8=ɯ�l�d۟�ꗷ?�����4��y��d�R2�ǥb��_�����'�k�xiu����VV���Õ�d_7�'b��C`vQ��Qp�]�z��>:����z�����С��K� ��y<�	8�Oŏڟ^�����K�X���b��x�7�³y�߷p���� ��i|J𷀠�.�q��E�}Q�HE��m�9 �s���#ӽ|��3�q��o�a�T�������\\�����h
�뜒H��\<f��6�N��զ��x��&�ʤX-#�O׽Wi^	��u�
��ܭ���j�L��a[�n���d�� q�ک�����H�?�^c�˰c�3��Z�����w��b��?�-�=ag��C���:��76���<�fx���_j�s޹� ~�_�S�B���~K}X����V��m�R�������NH�W���ໟ�6pi�l�~$д����3}�ueW�<�X���������� º#j��#�A��$��J	���xb<6C( �\U,tF�
� �R<g�i�/���^�'�^��rG2ۦ���� � W��(����?Z�u�V-�ZB��S��I��$��^� �\^kz>��C�<��ہ-g$�[0�7ʻ@�� ��_#���W?�E�hwQޤR����,� �խ6��,Շ��-�t)�uX�{٥�<��v�8����mGH�t�5�����)cO1"{f���I��V�)��{�|�:��qg{aj� �>�J�<)�ϵI�
h���|��+]Z[C)G�<��+�#�UO ����+�����������H�*���8�,3T.��=
g��]NYc�e����nzzⷼ�Դ�;+��y�r��j|��S�pN>Rq֬�O�Aԭo'��AeV��JVFNI�:�=s�.`8�$vh� Յ;�w�8��$�XL����aBǝ����Z���M�����$���6_*A
 �H�7$���֨	���6�Q�ȸ�1�����-��n��>?x�I�0}ɮ��?Mao.��\�%ݚ�r����G���=H�k��F�;]X�=��F�5S-�#�9,H�ԩ6쇡�k����j��olob�(�G�23�_Lx��
㿋n|0<;�]/P��d�����$J���7��̺��7��:h��m�V���.$M�2���=kꟊ_�O�o�/����#_��T��O�BrF��r@�`G�ҕTL6:��ڳ◊4o�y#�.�so���^��,��,�~�!Nd��^��۟�ŏ�o��t�N�\�K�X\]L���*�/�2nPz��{��K��NM'C��� �5�h���qI�h�ե̩��(�����<x�k��o�H�O�;�[}g�~-��ť��mn�� �(D��e9#����X������(����I+)���k�9c�$pO'�k�,~�2�������������?�]KDЕn'��{����`���B��T�C��*�7��0�ú������A9�ح,����q����� �����?	͟C�`?��u�?	n�P��t_�DR��㽹��~4h�X�=�
��ݏ���{��� ����7�D>	�P�dh�%y�&��8j6h����G������Od�I�1�����Rk+X֯��N�-m�x���d8޾�q�
�FOWc㚸��&�=�_d��˂v�^���J��	�Eo)����W�O� Z�5�au��u��]��,���:漋ǿ �q�mCJ�������{�Ĳ��NqҼ�V:�	)U���Z؍)��x^H��e�F�r3�����j�s���h
����\t�ۥqɫ���_�Ŵ� 4�xmx10�o�pk��|L�����m�]�,}��O#�����0��z3��aj����o4d�	I�P�Q�;�5GHԵ�B�;�869� ���[xєF�.ǐ+�RI���]	�kA��~�s����� l��?Z�g�^o�_�>x��������6V���+�N0���$��	<�W� ��y�x�uW�ԋ"n��6NnE|��<�l#�ぞ������x�|����>O�U϶��
��Z�N�� ����M3K�O����(���`pv�����⏃��y���h���bi,�圢�ɝ�r��+ӯ5��(ؖeC�H�A����ŁS>� @���W�)�">�� ��xfmkK���=:���q�ìM��K��UX��.y 3�י|����l�����>"s��Է�Ш6�ƈ3�  ����|��P���$s�lw8�5����������	a�L��5���S�\�錃��ԩ%����:ƨ~�跖�p̗p��碐����y��=%~�l��\Fc-���?νc���� �������isqo��c���LגOwy5�����#>m�%`��u�T��Z����n��$�e�H@*���b����Z]��t��ȲOi4����Lf��X������Vn����u~�4�KI�L����$.s��=뚦��rc*�$�E�;I R@������O-ăa)�x�Wm��p��n#�ĩ����%�X�r��=B9"ީ�L,:��z����o>	�em�����-����['̤��!��0ޫ}��ذ�Sin�$=��>:}sR��rN���#��}x��~fn�ұ��S�9F���&��8䈍��vJ�-�Q�����?�֒Y26� �W�&iW?2�N┖��ƴ�� x���o�D_nUzi�O���Ҿ��x�����6� �7'�uI�?�}B��^�;(����Nxm�G��-V���Җ�ƀ#|c�?ʾ0����H;}��_g�O��W�ߵw���� ���X��>o=� vG�j����9�q�X�"����c�%#h}�m9�?ϭl�J�M�Fr�~��\ιh[E�����<��8�yt�%�}���6��6�r�$���r~��W��c$�F=���h����#�9��+��?0��g��DU*���m��eQP,Q�g�jvO�����+y����m�޸��4���1��i֠��$��F�X308���-j��p����,r���n�����z#Jq�j�%��{J�a=�[8�+_��K��Xn>�3�ы�b%Hנ<�����n�P��V�kqC�2P��#קz��?k����[W�*=m#<O���r�����9R��~G�P�Q�*��o�?�޽�x�[��!]���kp�ev�d[��#)�=+۞�.kb����#��s����/ڟ�5���5y�q-�%���?�uZ6������Ś>��˛ �c����Q�{��W��,W��QG��ϲ軫���o�x�{�H�TףY�_cUTX�����|�c/�-g}mi���mJEW]2K�5�!�,����^}�~ҟ��Z�M�%kk�IZ)��ͅ��>�9�+����ŧ%vb8�y�_�����l+��8�j��n����<W���M�k�dh1�<��#��J��i?����~4ؿ�U�'�ɿ��\Q���}�5�˒[��إ}S1��q��E|e'�%��M����a� �*	�h_��$S�$��0�t����d%s�$��H�4��En)��)E&�G��?�k�mp�K`��=�ֻm�H�\���r4��.� U���KU�>Y�h,O?����(c��A�0{�ϧ�}����V�c��^ҫ��)>���<dsQ�2�6��f���h���$��{*�J�0?���g��b�a�ћ�� �&i���J�S�-��+����F���@��z��i%�����q\߆<�G�U�j�,���1�a�Dpy�
Ĭr�dp=j�ڑ�φ|T�g�ٗ���B�!��}��V����XW�R5~�q,���S�Fs�ʦ:�^
4��T���i⫽kX7��F�'��D�[�������Z��<aq|��~+�gh�1h�F��a������^Z<��:�9��Q���v��\i-�yU���r�����D�'��'x�Sa�c�Z�?�/�]L#p@�ڍ����U*	���#��;}J7�&	$\�v�
Ľ�u��8��}[��0����ݿ���]���"�^�kN?\��DK�;I�F��b��Q��?}G�\i9-�lN�U�q����1[yk�Y]��Q�}k���&��^Mi�	�x@�ő�ӭR־ Z<Zh�1�c��,e6��bh�)�2�Л��{O�� k~�5q�T��6����eޱ�lbrp��𪿴�Ŀj>�{�6�-o��D�� �%#����}�̼���?��N��&W���H����J��O�ڧ�_hv�xJ��K�LuI%W���o����^�0�5u�����N�G�h�a��o��Av�]��b����>���e��M��l�k;>��s��c�W�������7~�!_��j�j�8R�{�\�c��lqX;!H`AG��z�y��4cM�X򲼶�
NR��B���������#�O�FР�o�QɵT�5�} �6�(��C�� L#`Np1��	$�7d�<
�u	�M��è�Ԛ �M"��Υ�[�%���p��G����q[��sos0���1]���O�	ӭ�?�jSK���%��ߺـs�����XQ��_|?o=����o�)�K6�p6�X�q[��Y����@l�&���������|.�:�,t�Vm:��2er�$�J�C�\�sRh���ck6���-@6y�ȄF�b��I|�z|w��oss"�T�����Ͻm�� ��/�wß���X�8�k��:O���8���g��+�����<7�h���ֺ��J�+�-�p1�{�����'�`� ��ES=ƛxƻ�g89�2Nx�͍/m��w�{��G8�'�U�Ȉ�{��-�ŉ����~��ה�ci)��b�����1��s�zw�/k�ҵmj���z�cw�P��38b�%�(W9$��4� e�����uG����\��6��DKk��2��W�8*:W����5��,u� x��?ti$�[� �m.W��y"cX�%e$��sԏ~9]�n�>+���é
"H��ì9<��U�������v:�ϋ5�-rk� �Mg������}�$�O8�_�����T"+�[���D�gّ�q�1_����¯�֖W���<�o3ºz.�!B;,��e����y�f����G�m4� �c�ލ-܇N��G%�7W��4�wcp,s����/�_����15��t]"�Z:���Y{�����D�:��$@ � ��_��PҼI�íXk����������y�v�v��� ���J�6�� '�uT��o�������@�����_�C�τ5[i�������u�������$��)�d"|��z׻|n�Q���OO��?@�]#�1Og�y�E4/�2��e���W�x��rd���W�����j|^$�1��maI��P���*�4����d��c��k����_B��'O����T�� F9�k���O�)��'7��}b�v� ���N�Փb��6�ޝ���O��ĺ�^� �Ғ}�cY�C,�{�'ے�� s�3�J6 ��'[x��F��r3���P��-�}��۝÷�sOR�7��H)�p{�֭�sk�����Xٙ[i�R�X-��ݹ� d}j���M��>,[~Ͼ�}�ɢ�xn�F�.&�{���BHT�����#��Vn�7���&�L����z-7t�n��P�b��V�?�CcN28����h����T���k��ko�F%ki����=�) �A�ǀ>j���O�L��y�k�Ϛ�t����;)?9l������H�I�1G��w���RѼ�x�V� �TI1KG��.����p�wq��OJ��.%�a�����&y���Jd-�y'���ҿE�����{�B��9t���Mqqp.vRl�t��|�5�宽|<'):#LD-�o�n2���[S؉#F��@�<k.��=ٺ��&������� �F��<Y����Mfo��o���,o��x�z $�O<�8������,M}oix�en{����#h����L�m���u���t��[���S��prA���Ӑ��R�HM�6�ߗ`mm�ٮ`���?qK�ӷL�T��D�A�f�������O�Sb�9�_�ӵ_�y��zl6�-�i�z[B�'�I�����L�2鷑\E����"�GS����T����8�$2���<u ���4�#�f8���nQЁ�،֢�{V�M�P]�l�o�,{�޸��Vw�n�k{�!6��	3_�ts!ޭ��W��O}���uj�I:ܲ��T`,�����W�4������(m\���	#$�?�^ռa��s�_E<����	�ؤt�j����l�b��W��R��G�=�y�^u��h���N����J�`��n�n��B����/�.����`��K�4��6�v��H'$����<��ty�?h���twn��'���q_c~�������	��SY�P!-�;��Y���1R@ �����N��W"g4~*�4�#�u�{X�-^9��&�XH��א<����i+�'kլ� j��C]��A𵆕���D�f���ߖ`�NN�
���~�^�<�V�Q����z����4� ��%nq�N�������}Zh־��Ɉ��cA�,�̤r8�AϦ+	A[sD~�H�f���x�P��jn.�U׵r1w~��:6��p[��������i��!��'�L���gY����cP���9n̑�Q�[B�"0� �����k�uL6{���`�?ʺ���2�������6������m��M3+~ku�ƾp��|d�q(�I���{��B��>��҂�
�Do�C�1��x��Y��lM�8��'���5�l�����MQ�o�(,@�\�׉��n�Eaub�#��5ӕ�ĩ"�W��yZm?K����x�I	�}�� ��_�]��|��H�ḭ�:�Ա�K!�nq�Q�G<s����	���SSӷ\G$h�4<�@���p���{]��Y��;�+9���ƽ��Ŷ��d��ZhP�!_vy<�<b��+K���}�n�iҏ/R/�~1��+�����<�y]~����	�#�<�)��|g~�V�e�[\]\"���R}O���tK�]XbY�y}��[ᶯUf�䚫����Z�jV��|N���H����2ڳ��aovi��jї?c��Qh�Km=��u�����ݚ�,��*Λ>\���j�4_��q��g�x9Tg���s[j��
��=���d��|=��|��rh����l�+G}-��~"W��S�;�O�~�3L� �q�W�4Z$px���&�M^&;�3/��I�nm~���~�yi56}����Z���|��/�A�?|Z��M�mOE������s!f�0���P���[�#�H�'(�xT�b�'��%���ρ� ��?�c�M����]U��$�nۘ���^5������3�O���K���Z=�
�u	<ͅ���?�z|�'���F���3ѧ�K�F��M�Xx��Qh�L@�'�ǅo��$�W�x��X����"���*�x��mz��.�vV	Z$v,J�Ka@#9��忺z�涧�|W��J��<]�|+����J� �� ě˼"U ���1 �~P@�C�ſfM'��_�h�?j�ǃ��u��w�!�I"�2�ʩ$r�#?-{��/�??k������|g���>�7��E�1n,�sn���I�1^g�����_���d�s�ht���d�5�@ź�r	}��:�T�˩�a���>�$|j~r#�(����^��׽�A�R�mm��g ���q\��x_Y��Ʒ�ܪ��
z�؂+���֟7�͵�YQY][��F*���u~	�]�O�^"�E�ײ|ɘ��=�ԯ����<�n�c�x��~�V%hg�V��O!N޼ח�)����	�c�z%���?v^C =H c���R�g����7��N�|����v�:�G~O�=q\�����q��Ԏ���o�~��k>1О��ݞ巸Y�ub��{�Nk����Ğ��4��gym09�)x��K��?�;V�cKO�����YsN���/��j������S^x��l�HE�)���q��2J1�Ϟ��x�*����~�7�D�x�b���ǧJ�=���u~�>�h|����[;��.�;�NJ�����0��"Z"��eYFO~~���M�XkZS�����n@D����7M���Mf�N.���(���t3~̾; ��lQz�������sۏ�FTa�"���nM=mOIi���	C�l � �t�k��׵�k�xW*7	!�elgwJ䝜��1\<��=K�G�?|��ց���{}�N�Cj���pT��z�׮X~�~�����H�v���3c8������e�G��8x�]�t+[K����E�*�ET#9S�X׷�~Ξ����I��b�=�!� �F���L�{�Y{�q�A�;�A<o(���8��Ҷj���[i�E�bs���;~Uv�W�u� =)�)�H�*�{I����ڶ2���g�����}��?ʾ.���� �������a[Jl��� ��z��5i��H�?�w��{/��\���3#������]�?�⯈�F�嗉���1�,���=���m�|O�#ƚdO����H�YLn�d��^UIMw>*���u��Ǿ�]�1�v�Y���x$m��d�S��S���Ѯ9���0,W-��� ��蜩Ľ��(�~�9�|�3�e� H`�#Ң_�L��S*���I�T;KHv�Gb@ϰ�\q�3��|H�\q��q>'�{����B8�������i�� �iu\�����\C+H)	c8_�r0=����O�7S�<M�G����%�62���e�ː3ֺ�Ӓ�3Z�-U4�d�ϊ�u����4�}7K�U�)<��Px�cޙo�__[�宑uf�.c��Lp�!pO9Ǹ�C�~�o�[x�űͩ���#Mm̌P��ʀG�k��_���O��<0�zm�sb�-U7�1��rF8����g�O���4�Q�r�~�|��:[i���ċV�޺<����ޣ�]T�/�߃^=�Z�Euo�X��a�ܩ8<��v����x�o�vP,�ʷ:lq�I*9�9]�6�>����z�ޔ�}�B���0�G����R:�jף�YT�� �H��]T߳O��K�r�g%��g.��x��o�|m{w�OIS[h�U��v��Y�U*��Ҽ��ڶ�y�N�X��J�n�2������v���^M}�O�4��>,��a�n-l����9bO� K#����۴��9C.����%h|o��ZGus�^Z�w*����dL�¶s���1�N4��;�;^�4��G˳j�y�p��-���gI��5��N�������;�}s�f����[���SQ������f��uw#�w���}+����H�kڠ�S�B���4Kx�[��K1]��c mǽg����r�g���`�g��畹O�f���[��ӯ�8k{�?�?�$��i�ǌ��#ھ�Э5�|-�n<Eq�-�4�����h��̡���Np�ݒ"�������7:-�ƥ�qK�\���ʿ�-f�Lw�SJ�Br�����,�!����{�����\|��BH�=k�񷌓���f�D����H�",� ���[Y�����i:��Ȼ��m�7@�n����]�#GO�Z5���L�%�g��V���\��z}+УE�RG��Rz����/�vi�k6��Z�����TH0z���=��z}އ���JA���KL���K�t鬋�Ж H��X�c��5�������L|�:ͰZF<����V�爼h5��5K�zXZ4H���$�;=8�u�6R�N-v�.��j��zD�L��0�T��P g$������ֵ[���2R˼��s�?���u��+�M:9�Q���������28�f��h-�b�M7�4Y�����#��n;=Y��r�l�4���ûM[N��':��@/�n�y;f����zׇF��kWV�� �0En&]��S��Gę
�.������Wi������
G���Ǌ�T�-�s��:iX�o������k
�mH#�8$�>n>��Gý×�ڶ��5{�kD]���0X�����
9<��N���vg�e���}a^su��.)u;8�}�S�Q:炻�r��z�5�d*u���7��G���|	f�i�1� ��G��v��� �� �֫�������Do��x�I-u4�rOP	8�[�ڃ��-�Ķ�$� ���a_�I	���<���O�x�N���h�Dv2Cr"*��n��I�� �W*n.�c�N�oS���_Yey�5��+g�tq�-Z�|:�xn�m$Z����	[yf*HpI=28�U�x� IӬ� �u}\Yj�̮��ʏl�Һ�x���t��H��`���Ѯ@_9B�Tu5�-��#��&��ˡ�5ɻ��gg2	\� g���W�t�>��,���]���YI߽Mi�� ��O��E�g�u?�4���t��2ێ>q��<�y�ܯ�fo��I<�i0�y���Ё������W�N��G�4�(х��.!k9�uF�vH��A8�>�o�`HY?2�֤�῎�� ķ�~��3��i���͟�S�VE׈-,���a��I�$VS�r��n���7����9$�d
8�,z
g�#%�y�x�Y��7�U�3��ua� }R/��T�!@FpMW4{��� 2.H�æGQ���-�B=��lO����q���� 	&�"�I�[+gj��Ar��ŅӺ�y����ގd_���3�|�Kx7����76�텓_>�$��6����z� �J�� #�ma��Ē��S��������GJ����������h�C��%�������x����V�[�;��]Γs4BhDВ�F�0de�#�r�^2�L���t�k���O��qu&�.� �P����8�*�dq����<��Nx �"���H���}JL�_��S��G� ��4/���[�ѭ���idl]-����c�v$u��q�#d��+�Ϫ~����%�0Yt��|���Q���p�q޿6��'�v�cc���/�[{K;Rdy$s��=�W���/�ؿ⾑ugqo-��y!a�1���3_�?�$���Io�?�r�f�wfA��8���+I3(�w���?�4��|1ն.:O�2��F1Mo�7���F�Uda��1�$��)�٨�e�7���W�_!�Ŧ�acqm��j�β#���v`�V�^+�!�� ���~=�c��hZN�o�ȧ�0���C�ʏZ�ٺ���U���6iĚ-��_I�$k1��ɧ
7 �>�������<5�X[|'����ɖK�[��<�y­��!G'�Z����㫿h�;���>ݣ�vMF�;�tYF�{�{~�7�?l^-/D�ڿֵ�f����F��+��*�%���i�9����&�����FMcZ�4_��,��{]�%�֎�ؔV}�˖c����z�<!�[�_���ῇ�#�t�,���M�X�)��m$g�k�7�]���k�8�׋.�ui�e�����X<0NM�d]��8!���\�<)�xJ�H�=��e�֮��T�N[ōZ��m�PĐ��QIJ�w��m�/�n�Wx����G�Y���N��9>��>$��/�z�߉<��4	o�4�,�Ws�3�OL{����k{����#Őjv� "_YyQ�1�
�T�g��z�u������ �'_ů�r�K�[&�`��$�7O-��*÷�Թ��?.���ĚZ�Z�u�[O�*��Zd�����uBpj��)�J���o'�$���ҿQ� e��w����ÚƗ�}N�y-�SԬ��ƪ�D���0��?ÿ>+���e�º��-B�E>S}��%>Z�>�g���Z�~Sk�|g�;�k�״;���:XS��,�g޹y�w��M˸Nz����5��㯉ڗ���&׏�I�7���^��)d�<���:�0�#���_�K5��Q�5P]1���}�Wv��>���˭���\�MQ|��3__��Fn��!0��8���ރ5�^)��#�}B84���^u��1�ݧ�G�f�W���'������ ��G��g�kOhSO���N���v{I >UW�c�0�2O=EG����n��o5���-�@.t����&K�(bE��mʒ�8��$���|Y���ƿc�{-V�|!q3�u��<�-w9�"��-�(���/$O۴(f��D$����_t�#�
��Yh�o�d�%��$���� ԕ���]�p��~A�_x�ƒ|Fկu�l�SM.�]g8<���tA�c+w4�=u�Z��wce/�q���	���	9�lU�K�=��۝=�YS�7�>F��`q����?F����5�ͨK$�WO5�biax�Pr÷��#�%�tټ��{�7nf�>�cWBĨ8 �J��2�ĺ曢6�mq"�I8�;��y�Ƣ���V�uBMB�h-�,�I;�0	��������m�h����Eq���:���Z�=�����Y�v�e0F�iѠ)%NCE�E��V��I�i�֪V��^9�S������a}}6���qi��Y�y����/���靾����ȴ�{[�[{��E�DDM
d���G98�����s��onb�b}�[�D�{��j����YY/���Z�Q*�%Ě�2H��B~_ֲ��+{MZ���0�mZ_4[�H(����5�ɧ$�k�M������vJ& XnI���+��i�+c-�V2y`�Aц}r{�����Z��#H������!�f�� N��^i6���h��ԗ�i��V�e�ZNATFO�6:�W�\T6>(�����Ă�o%��n>��Q'�����k꿌� �Q-?�W�H|9o�sg�.�bp��ѪK~�b�3��ѲzR�+� y���3�x��M��t]S@�̖��_Y��ǘ�x�Н�2��{|��N/ȷS��#Դ�?s�5̾!7
�w� �w9m��I�������<)�]2���~kV?����f�BB��\ݱ�`�v���9[�I��/�	�E��YA�����||��į�$q�9�}��#������R�5oi����[h#c��!�qY+���q^�\5����q�Gs�����7�'���MG^���V������M�+1$nl�^=����k)����j��we�ۛ[�C[�m�!���=;b��������,m�g�	��L���d)v�8_��8�_4���� ��.�� v�1��./��IYR_LLc��ŏ�����l���+0��a��L�5�l|Fq�V;�oRx`T�X�}6�IU\��\��N�W�|=�Ɓ5�R-=�I1G��f�$�A r*��k�o�w�jV����-���OE'�=A���#��*����|��+s5������I�4�Yo&��n9s����k�xN�oR�+eiaFXez{�6����Vi����/�_ֱ|W���tMb+��(�I"[Y�r����8�b�}b��{�K��=�8Ӫ�9o���V���K��O�B�����V�?m�u�5�B{�e��ٙP6pr��)��G��"��h�|��f3���e==���Y{���9�w�s�n�p���)ΎTUk������)-��xD]��L��yܽ��A�[��b0Lc���V���=2��'�Y1�v�\��@�+6�9� 8��G�F6����|'�5e��R�#�|�-�D��\�N�}q�G'�}e�q_�~�������� �y@c�s�?`�|w�z�6���'��9$�;[�d�8;IpF99$+��&� ~g�9;� dG΋f�\e��I9 a{�� ��o�a�g�zQ�/<���E�G��	����� ���{�Zo��=���� �m�Aim��������q�5/�O�;����S��ea�]&�Z�Z�� ���2>o�j�T{I�#�XAo# �Y�%�q�~޵���?Ð��&��c<��ǆZe$�3��O�⸿��?�� ����K�Ke���<���3�"m�����^�� ��H��m�.n���0G\;� ��� ���s����W����'���4)w34M��/�eF~�Wi5����\i��M��B�5둎@q�W3��dئ����P\o*���:�� z�Gk�"��{�nf�|�P��8��J&4#Ie(���$��(��:z�j�~ɭK�l�\�y0�����ߕU���4��G$���@�O���+A�ׇu�h쌇Ov��o3<������>Tsb�9В��λ���σ�.���#���.c��9�=y���{�qo2�h�f~rzs�fj�t,�Ym �fa���G�
�][Q��X^X�ɧ���t�a��kş���+`��O�-�z�kMt#V��op}j^y�k����یsX��rӉ�l1�co�qߎ�i&kƸ-����s�ˡ�:5a��6_�|�t�v���|� ���$l�m����"�O���]6��a�M����<@��x��-��l�,n��ߖ�s���T���g���O�� �jK� �G_RFr�������$�#����=NBc�J6Qz⾡��2�:��n�N(��&����d�,�L�=F9�*�{c�V��)�H�)OJF�@��R��� *��������~���_hHx?C���ڦ)f���[�Ir���j��5s�%�I�����.Xt��G+��Ě7��][P��.�����Y��np���z�c�Z~��B�Ɵ|G�x�]�MI��,�#�Ь�\*잸#q�\�Ǆ~$�U�:�o ���'�2H#�j�u�|P��Z)|9��I������kå�тQ����4q��$i;2��3� ��%X,�y8����|��M.�S��SO�����#X���x�fy#�Ѱp�<�n���>g���A�1!�	�YVu%]3��P�GJ���)$�H�
�]]��<����O {� T�1;(���|�[�C<�x̍� �޸�ӽe�L�Ni=�W��o~���g�+X���Z�"���	F*H��W=��<y�<|6��I��=~i�[�]cVe�9a��W��_��-ʾ�t�9.��[���p�`���c>��x���/����:>�!XR;x,��0e7�I�NUaF;���֣��!�����i��
.4�c��VL�I�W'�n��2|b�<�V�c��6]�|�N�o�d\�g�G��+�5_�> ���� �~-�շ�n�i�u�C�gU� #��\-��?|P�������Y��\_]iۣ��]���� >�1���$}N�l����oX|B�Qg{���x��Q4��<��o���n6���)�����};S�`[�t�^�+��;�w��s�?��H��+��~��\�6�L��]8� ���{09�.05��_��.�y𾠺���A�XZ:����H�>Ƹ��x�2�>�t1��hԎ��/�����@��� gLHیeI����Z�	g_�q�6����g?"����A�
�?jO�H�?��ڣI����䷒���9%�A(W8��N9�5��#�K�h�
�Ox��a�-�nBfr@����X[���>��XnW'.�C�_O�x�\��f};F�{�uݑ��#�O �,Oz�~&��Ꮛ��4ˁ���� �~A�g��S�_�p\xJ��R�����=�^���-��8U�lgk������7��{H���i�#���ɔX���d+�H�y ��C5ʱT���ݏ7.�)S��SK�{�(d�ោG�c:m��S�������5�-#��I(T��Ak��<�T�s�s�ִn>-Z|)�7�-Qu/˧���i���� � >޵KM�{�柣����gV�]�-L�J���1�������Zuj՛�93�f�S�1���R��h������-�Z���I�{e�0u�x�\� :��7�F� ��ň<R�7�n�[����Hӄ�k|�䃁�9��/Ɵ<|���������r���.��c`������\���-o��~#G&���VP�=��`�U�H���cvy�x���7EI4|kB6Q��<;�&��s^׬g]Vk�#�|=;%��B�^@�8�=���� 	Ɩ��>1Դ	��m�-�J�x`?�֩�,�k?�hw���:N�d�
��c��c�j�x|E��X��K@��n�������9��r�);��,D�<���BMb�N�f��K��^��B`��P���U�8����j���ڄ�r�<�;N>Q� ��k���xL�)���T��6�bڧ$��n��x�J���/�RO68\*> ,8 ��5�JQ�G�RN^�Cg�+���-����k����)����?����t��3��[���k�қ��tm���Ӛ��i��Q��v��#F�K9�"��څ���7����\�#,N}ɬ� x�O��{s����F�J��Z��>k�t��!�-J�<�-X���z.v��tT��M��::s&T��m5���H.n\	Y���9�.ߕg���S���)c��q��j����w;˻��ד]������}�
�YC,��� }�� ��ls_�?�xW���k�Q��v�yRk*��Ȍ����zױ��)+7���~O,J�Ilxw���>�o��{��mGGFk-�p�#dI'�N���_��%����6��(�u��o�&�+<��㟓8�}�U_���w�~	êC6������;+2���n��'�¿"���>>��N�v��J�J��w�\� Z�!EY�P�Ӥ�l}�k�
/��WRY�F���d���@Ӣt9��J�{�����)t�G�F�=��m��C�M��3�j�c��S$�\����S�Un�H��$�+E���k4l�>��5���i�8֣�J�f����V
ą`��1��˞��h��'��:ݭ5�;�:{(W��=�w,�y��`H��$��&���B0���8�V|�mu�^���׭1�rQj�]Bh�~x����s��Rs��9g��w��"���Y�7�.|?km��m��h�9�6�i���s�c����J��hD����s���|8��⿄m-��r5�ȯ{�_�Wezn�pB��s�iю��q]*��L�.�4��|�-��jX���g��1&��o�z�����5��q�o�=ލ�]�>�w�^�h��g1?pJ挒N��'$�>$���ӥ�V�G�m#(�3�� ���\ן(�2�gϪ5p�Tdϥ?mKx��^�f���G{gq��у�q�s�zW�����_��G�4/���x��� U[�-�@�Ф�A<�P��+�?iMI<E��;V��b�%�dg�Si+�=�A_G ۝�GNG�=+ե~]O��� w�$���X��[J�BH\}�O��'v@���O�Ҫ���W_5��� jW�v��J��?���s��V<6@ � ���owm��� b��-�D{�����p~��}�����ݿ�-xCX��-&�M�-���.M�dd�o��~��+�׌g�m��x����A���-�*IC���#!q��k��c:F�"]#f5��p0;� Z������3����I���f�!��?q�L��Lh҉Y�*�['�4�dz_���j/�|i�Y���Ο�����F������V�31l 8�_[�I�<k�]z=^����1U�#K O,7� ��8"�Y��� gM_�v���
hz��O�7�m=ޘ"���w�z���8��Ҿ����K='�7�n��&k_ �H�w�J;�8#�#��o����φ�2�M<��|C�ޝ�������l5��Xn%>b��8VA�x%I���� �����M�'�g���#�˽��)�1�+H��c�N�,y�?��� ��]����Z�t] i�]R}OҒ�+�cݸ*F�SzG��9l�sK���<1��M�4��Z��aq�Op<�o0VV��p�yc�t���c��g�� �_����/�o�����Ok�ic6���[�-�,���H8��8�=�/�eo���Uo!�n/����6�j�4��,y�y��C�����.M�;��-��h�Rx{L�p��~ޏ2���!���#��5�� a�J�Ꮔ~"Xx��>#���-ti,��ʑ�� �
�<��sCR[W�>����|I�� ��|8��.,m��_j��	��1��8��G�u�x?�a���N=�Q}n�f��,�DK+)e`�)C��8��}M�|-����ң���\$Vе����͒�,��8��f0@�s��;k_fO�c�����n��6�K����h�ِ)r��j��u��h�x��W����_�^�B<=u����RO%��>�<DN�(�}ĸR6�����ݮ~?j�uO|-����b���"nⅈ�[�8��ھs�3�x�X�[���:Eƕ�7�����Љ���x�,T;�Xr8�:��>5�7�;�	çh��<;s%ݻ�u�hQ�Z�l�-�Gk����94�.���8���>�0���e�{ᾧ� 	~�⻙���le4��#��eV(Jdd�����)eas�&��xL_n��-�i7�럧�/�[x��v��g�u��h�Ş����#%�R*��v��v�7�����㕣���WS��Aܤ�cpx���ϡ�å~�:F��f��^�|Q�YE-��E�ܠn�%��6��|��+�+��
��xk���N�~�$cQ���T��rNO*5I�l����.��-gV[mFI"/|�-��2�Ѱ+&�6���n=�?�_�.����u_��P6��z�I��g>��&Đ��<6���l� S@��$���G��G�	g�GC�<E�����p����=�20�n"�7r� ���Z��5?��N�F�)J��>�q��mv��k�i��Io�Gu����X�1�5�;wE�ʱS���	"�?T�|L���w5��6��8=��{ޚv3��~���oæ����o+�Ť��&�
b7t��c��ֺO���t�5	��M��x�?/ha��Ϲ9��:坆��Y�ir��g)�)#�G�l���DTz����Guw�qcy+�%�5oM�G\�4�X"ޭl/��������3琨� 3��1��_i�j~�޳s~��Cr�G2��bP@Cߜ�}�i���b�:u����H��� �	!�*py�����,*������-5ԹI0,�}��K�cM|NH~ߤj��n5�`N�$c����I ��ʹ�*A��Z�Ưw�ꏨ^�=�R5D `*����6��ʼ~�r{V�VD3oA�қN���]9��u���"��� ?Z��V���Q�H���A�u=ww����f���>j����l�Z̪�1����CX�#�5F�%�8���tFS� �v����C��º���9i�#}CU�"������g�����q��S�3�ՓY��ω4��D�b��X䈱�V
�[���q����}��� 4�kL��Ͻ�� ��.�#v������^ ��~-|H�����\Y[��%���C9�
�q����Np>QԺ���GT{���f�x��<�-`���$�d���ː4��V�#�U,c��$���k�8�ƥ{���3�0�
�uw��5�2��xÃ����A���;�� ͤWĞ9�����&;;�%t�-�6�e{�}�ی��d�<�ƛ�v�x��7Yx_�r\O�[�?�P3��`nC.��}�s�W<�KEY�0~��><�7��+�x���Z�l�I��Gm5�+��%ʄ ���� .N������؍Fu��g�\oEf��.�I<�W��w��~,�����氷�2���	�"򪓅�^z���W�/�$��t�9 ��%�Q�/*Xt�?馴"[3�����4����Z�[�xn��[T`��x�t��^� �O�"Xq!�(ш\|�~��_@|v{m��mm�Xn4k�V0��R8�����5���x����-����  �J�'����|^q��ȏ��υ>6���>��柨�Ei,;T�ZH��7�pz~���k;�7[���<5.��ɨ��/�i�.#���u0��K�D���oa ��;�sC��l���)9`�3�����Q���5_�_��K9�T"�[{U�~ؤn�� ��O�4�xc�Я�ɵ�\�����[oE��"A� 9�=S@�ba��wc��ֽ�%s��m�>]=-�I�����VÜ�zT7�Q=��$���m�������ф�2�DI;L��i�~�$r'����$�'Oz�%!�4���W�X'�ʄi[������~���F�{��>ÿ֖�U��b��T\|����S4w��S�x�y����`}*�U�ݚ<��� �<#n�*5��{�@��ת��T��.�~+|�<q�����xbp�O��,�_d�q\������>�Wɒ���,ja:��z�?��_ş�zƉ��-��q+Ll/-#��1�̋ ;wq�zc������?K���$Oү��`�i��ޱ��
k^
�m3�:���ͥ�4�m���$�s��	���x��?~,�x�K�����T�D�a��;��H�/��� m���?���� 	ZK�=��q�KH�� ���h�r0y��Z���q�m�ɦA�k~'��O�t�d��V���C(vS�\� 	8����]�VQrV?J5
�_�Wᯆ����^5���+{�$��1��|�y����9����Z?�?�Y�XZEa�R̖����]�s��ň��k�M���Y����x�I�oj�I���,m�b c�O'?M��~&�~*x����G��6��<��BB���� �:UE�J�yc��f��u�I��
����[�?����|�2X4�֑�� f#i�yy5�xWO�=;Z�SP���.�C̮A�>���^��-�7o"O����^j�=����h�ٞo���&�0E��o�"WN�����$���6�J���7��ˈ�U8�����՞�߻/G'�Id���/_�kV�.�'�� z�*Ż��8���^}xk�}ԍ9K���� /���I<U�gO�������گ��G�r�rJ<a���E�%Nx�j���K��E��̂ٛ�,�r�3���:O���W�*�36Ts�k�O٥�|����i��q�����w��B���$j��8��w��?!T�2hE�ryֿ8��� =�THT�l95���ھ��I��R�Hy�Ҕ��.ǝ��S�����O���h�Ѽo����|Ź���l�B���c����L[r��]%ߍ���c9����_��!n-��TV��U-o�f�H�=�r�R[�����gz(���>(���k+��L|�he�`�������'j���5�Cv��Fs�9�� � ���7x�q� Y���ˎ������<���M���1���[Z�#�����Ҋ_K4�2*�<��zWb�+�6c�Ҝ3]\�M��Zi�SH�%������k��N��.�]�I�브W�$g��i���B���X�9[��!����5��I�g~Ǜ����~�赩����s&�Tm-�*�����n��Z�����i`nLg��G�6��ѥ������1Y�+��Q�Z\irD��!�1��u��Ȱ�N��^����S�Z�eN0�����},~���R{��Wp�F1^7�}*'I�u�hX�{g�ʽS��o3C��;�S�>Q���\�v����D��}M}FCy`9�s��.vƾTAp]fe#�{����O�����5-�b�}�ݕ��Σ���|?��Yj��3��w�x�����'o��P��;
���[�R�?���O��x�`�ϒ�m�{�5�5�����9c��>ǹ���=#�^񽞙������9�T'��t#������_j�K�]xSH�uIt�i���Jz���*2z�5�� k-{���ѭt�:kkX���`��{�5e� m/�h:T��p����_-���ө5�;��qY5:U���c����?�6mk�^��e�m��f����%]�@��Λ�wⅇ�>� �Ǜÿj��uY�wi٦(I <�~lc1_;|L������mR�l�mD�1��0)��<�zׂ��i��k7͂ܶ?�?�}.[S�g,BI�~#C�Ia6H�_�+��Y���6>'�\�{��'���CF�N{����+o�"�}OH�l���H�QԘ	�� uU�e�ƾ<�i�;��"kk��U��.����t�+��z瑃]��9��╿��u������o2��I.�~f��z��F���� jQT��}��/�~��i�x����<A�i�t���Cr��W$�'F3�$ח�+���~��-�>+^�/���_�P�!�I��_j��K���d��g��ahS������}��|3��T�K��g��;h��#����q���R1��pc�b��R�Y��5����M�u�>������M���Z�� jڥ��KnO�*���S�:���Z�WԼO��kE��y'�~� z
�o�c��Z�Xi
8�R�W���m��r�i�DYO��v������O<���l޻�3��)�-=6�� ��>�.4_�RY^�K�f�y�Ua�=�OCU��7���.�������O�_l�����2M#���I�>���E)q��t*��oƾ�\�Q��_����7����KK������\Ʒ�t��`0@$�S��*��P�<Ew�B�Mmi�����_l��t���X���Mgxju�^� N���ͬ�]�"�ҥs�#��N�cЊ�ihg\K7��X��]@ڷ�����a�N5�w.�w=�ͺY-�����5g�5/f�F� US¨��Ga���ׄybx���dn�˻�o�O��� �vG�����t=9�O^��]��yS� Z��[x3º4�B�W��)�|u>��V���z�W���M����h�PIsy��?��~0��[�	�o����:7�u���żф���q�S<��W)g������� H�[%s<�p@�Qp>n3�2>������;߆���w��&GӖX�y0w|ܩ`J�)�mF=�k-��bj/e��^�� f�M��0B/&�d��s��#&I��8�ۥ|�]~����<C��[�Z��z�"�գ�r\�Yc��L�S�]?���X��[�v�z��f[�n�3�G��99�|sھC��,�2C����z�c]��S�b�5�9�={����`6��X�&����г N���i��
Y�r�/ό����5��>UYs��21���m{h��g/��FvYS'U���Msz´��K&J��ʷ���*I�p�y%���;�rZ�jBs����Uǐk
cތ0��W�=ktk�\0a���w���Z;���c�y�s��.c������:��%�v`B��qګl����n�]]���EDߕ'(��=x����RG�"(_S�=Dy�O.�p��y��q�H�}A�G��kּU���r� ]���g�n��o:���%��'n2G8��M[N6���\� ��fZޮ�t�d�q�J�O�c�Ǟ�'Z�pS��5l<k��s��\���N�?{%� t��Ҿ/�m���ɯ�ڃBM�	����k�x��ʸT���A������%�Rx�Ȫ��F�%5�WTdS�1�F��SK���w���������|-=����It�:��Ci�ĕV$�8�h2���[������u�\�8{K��it�9
͵��# �_�߳��S@������\x����O�b��y����e�
8�w+:��˟���?��T�4�h%�Ӕ�=��s$�!��Tx�p��ڬ|=� �d|r�4�Y\h~��4��������4o���lr0Iw��\����?�_� x��>�S����Q�j��� ��R��烏s\���O���6��S�v�In�����ʲ7���b@���zWƗ���<!�o��Z���#M���ү����X�1��G*cı��pCgk��s�w�������'ōkI��{�m���L�ʁ���s�0F*T��p3Y�/������SP��!��Iq5���-�m�;�lJfX.x�8��<)�?�W����>$Gw{6ɩA�p�� z`t v�b��K��>ˬx���͍L�I}yp�XSsl%�d�X��nC�8�ڞ$������Y�=�̶�K"?!N�����9�m_rb����xkǿ�[�M^��ZҬ��!w�#m�H���ּ��y��o�'� �4�2��X�$��B�H�H��,��`0��<�q�׏��*~ѿ���_k���<G�j6����[���@w$�~dpwC� p_� iߋ� 	t4Ѽ+��OLҕ�E�%&��I"��rzw�1���ϻt��㎏�N��Σ�Z۴Mqkg5�_�0��<q3)X������A�_�|!� �s|[�u�2m*�`�.��戀����z}k���p~��ݾ(��r�V��1�b�X�/���3�� �����-[R��eś�*ʽJ�UW?ÚT��7s����U�| ��,u��yq*���I-C�����g�p3K����eu�� kk>"��3ʺ�,./]�`-���F������k���� ���_�~�����kq�h6d�l$���#�r�|�o�q'8ɮ���\�� �P�?&�f9=G0��Ê�F�
-j���X�G� ����j�}$W�}��TM��EF�9�{�_��m�Z��lf����Xc��m��,��y�9����> ~�_>(�R��)��Ρ�� �6�1y�9�2($~5�W1��C7����O,��9�}x杴�u��Ǽm+M���� ��P�,�?s�Ekݢ,�Ң 6RT�S�_0|j���gx<?a{o�b��Fie��z���#���@�0zW ��/�� |��:ƙ�k;t�Վ�}m���m<�މ�����������X꒭ƕ*���,.\H��,��P7�H ��|�Դ���?�y�6\|/�o'�$��Mv]j���2� �;���&�t�\�,�;��i�H|��@��$g#�0J��M6� P�|5�K���Ѯ.��ز�W��W��#�xd�t��+J��p8�q��ޚ�!���ʰ��S���:Tp�c�7F$G�3�V.���e8�<�!���m,Q���W�޵$���Ƅo���2)�����;y?Β(�#*4�w�K��O�J�c`��T�f���4 ���Ɇ�ݮy�4��G��n���\Z��c�1d��ޟ���?+���Pt�J�2��1��u%f
a�f��#�#�q�>���,������G�k#�԰��R�_2\H���>���t>��~����^5��q}3],�q��,A�k�_��7�-��ᾗ�
x�QҮ&�Mm���܆ݗ*9'o�q�J�+�����a@�1�-�#g'9�5���zxf�����D��T����_��%�|Ȗ�	�,n'�;y��EH��⎇�z'�߅��A�w�� c�o]Gm�����i�+Dĥ�Q�2T/��B�WԞ ��O�iڏÿ�����TU ���#.r�������W��3^�<+���?�J\\�����n"2'����[8'?.q��<o����<3�d���5��+�k��m5�B�00�b��F6�=�\��~��։��Ưq��k^��./�f����pcP_��'\�~��[���O[{���yro���3��0�͞G�l�@o[����r\��i����>Y
�@Q��9�c��\�jҫ.[�� ���鄕��g���S��?,��x�V�t��~�ˁ��M�H�ȭ��+^i�/|����^��t���Jd0�h�H��#���k�MA��v�H���� |1�ě;��hw�R�ǐɘ�C��# �Fk������3���"<����c��[�_�����M���F��F�>�z*�Z��]"}��9��A��$<�l�#�l:�ɶ߲?�O\:4��M��U�.�s�q�ga���s^m}�j~׵=�?/R���M���U�7ur�<���Ã���5�ˈ3�8� �p����z?�� ����O��!\j��1� ���v}���?69�/�O���P������}d��:��捄�H(T!!��|��� ����x��W	�II{5�*%��$�2Cs9��8#��*kx��O��9xoX���E��#��k����Oq�� 'O3�b�
sH�鑖�y��]J�W���O�$���=������u��0 �H��a#���5��|b����~�|�
�<1r�Mد��uԡ�ӡ�[�|�o�>I�]G^��vZ����i�[�w�Ţ[�o���B@;�jc��`��ֱϳ��,����:W�O��3���^��i?�~���ي�5��||�C�hs_h���5u`#ҟCk]��d��`t�5�,��<o������Y��X��+�rɾ6�n���r9R;Wi���#g"�M�����m)�g �ⵗfMT#�%�N����˿��i��94{-<9��ߗ8����뉴��Ri[M���T�ֱ;�� {�'�A2�d+/��=5���"��� ���m> ��NX\�~ �����.#��Wf@�x�D�UJ��֥N8zJ�5��V&���KH��F
������	�*]J�R��Q�i��p�����H}p�+���W������x��V�Ꮘ�i�}N��\[�n$b'���U�v����R �ʖ��Q�� h�Ҽ���{�\�'Gլ�h����Ώ�����GQ�r�{�[ܫAǳ/?�}u� �6z��ۄP/LX���Oo��X��R�K;���p���s���[�f �1�<b�?��6�Ka���ǅ�#r0N󎵤�S�>T�{�M.���Q:�q,	�F�����O\�zv��]kK�m
�?Pc�$`����z�? ۼ�w���T�H ���^�aa�60]�����d��䑌�T�ܣ�x^��W3Ĝcj̄� :�~��4=B�E�,��ɣup2q����������I��W�t����~�"���� �^�+¯a�k?5��a:Eod����k���(�6El?�����$1x�SP��� ���@���ú\j���}�~�_
.&��o5O�m$�^EHr ��j�~Z�k��Y��Qӡ��X%�˴��Ђ��E�1��u2J�-�g�?�R-6��瞦��3����5�o�o�}+���"�>�r0Ol�P�;�mt̖��$�Ծ����@vu���)]V+�1U&���e��9$q�w ���2��z�,�a�Oz�6��7��M�nm�Z����qm=�)�`NC�*(|ൺ�(>O4n�f`�������M�xWgU�� � q� 
z���Փ' ��*���>��߂�{�|3��4_x!4�9'��~�A�I;��������ĸ�M����nO\�>���V�����,��hғ�G�j���}p� 
��[Z��Ϭ\-��NTH��ݪ@���]�����N�:�����z�W�ߵ��dҼI�H��s������_Ub�^��4[G��A�����$�1�A�>����+G���s������GI��,5��ũiQ��L�������~�c�+c���xR4-�r���1(+�dg�^m��������!4kX��k�œj��!���9���^<�#���8t�FX㑀$m�An��W�U�p܊���S3�pt״w���-����+��j��@�UtR-�-���c�1P|I�5׋�Y/�!���@�n�<�3�>�� *��o���֡m�����i�;#�2y'�~5���|���>SR�i�i�#R�C���翷�ϳ���2����$6�Cw�wm<�?Z�&��uf�f��M��N�H�p� ~H����y��������?X�U%de%�p��Ą秽y�q�l\\hO��W�k���^60�� (s�����1|] <%>n��Y�3h�H�+
��c���9��K�7K��֎�P��� ���Q��k��^�2n����W+Q���_~��_��B�J��/��,�īw�ǯ�]��3πdo��.����_xw�~6ԭ�B�5[�s�&�9<��p??:��~("�tn�HX�� ��f��ϓ�g�<ƅ<4c,���=�����-'��y�iQ��3�C�F2C)<��֗�1���e���	��Sl��1�O�_?�G��7P\x��S��ᶲ�
����<��~8_�J?b]:]5�h�Rh��9�\��e4gB��:���y؊Я��5O�����T��|!�(5�����IX�>����ƣ�u)5�VWJ$����������xKħŚL���A~�h��� r��W�i�����f�A$38��r���oz�U�	F�-���Zl}3�:�b�Gŉa�� �"�*H��^5�6xgE����ō��Q�$+�^k�� e[x�E�����:[���v�d� G�<t��Ȗ��!ׅ����ژ|D ��猫���<�s�}��
q�9�c�)?g��[�� �#f1���N3����r�n�'��;!�L�*����:���f�s�EI؞"�̎A�EI� 
��dv�͠��F�]��'�0s�9���,��d���ϧ��ѕ9/�=���2�@��}ea#Igk=�v�H�	���=�ޖ�s�xi�l�7��w@�r ����mr�P��C=�nx'��ã�Nw�VzN���GL�/u6n�["m2S���;s�J�ƽ�"�����V&R�W.����|=u"�&�w"_G��	c�WӐs�QxoH�о!]E"���n�V`W#��+��K�u�i��R(V�� `�a���gߥR�;Cg�ǣ	z`��F�=Gp�����7���,[y-�E"�>[�*L�3���z.����i��h�Ĩ��>#�cB����:�L3I��t$20�R�#�{4k)�������[�@� �W���s� Z��<o��)�#*}ԒA�+G^�>�w�ټ����[A�ſ4�w浸�>a��}�+�ST���g��#G�� ��_�4���&�5ER�
��d��r�5�� ��A��/��<�.T%��e�ŷ�R���F:�־f��t�z=wŋ
A��
�Iq�#1*�	<c�5��g�4�~ ���]?Uե�O�L�L��\�}�^�ʯn~���#J��-���n��%�/5]Bf�������C�f'��W�h�H�)9A�w����`xR�}���,���x�W^�Q_a\��X�^���]��V�;w��:-S��8����^����y�5VY�Y��.NӜ�e	sw��,��|�W�+*Yq��?7#���Nd�H�U7�$�Y�Qǯ4�n-af.����Oj~���S^Ho�d��E#��Ž���Sϯ�W-m�g/��{1N[X�Fm���n*����q��.������� ��:��k�[��5Yo?� ��p\�`V�:���%`X��0��S�|y��� �����H�^?�c���x��"���Ǘwo7�#�ǖ�Z�*T���� �sAH����]� �/�I!y$��of���"��k�3�u������>:�H� ��� ��ʹ� �N�� �U2�F=|kn[���*�a-��Gj���	K7�b���u����!�=8�?J���3�<����wƟ~�_���������BH����e�� �{֤���EѼ�� ����v/�Nm<;���G)��\
[b� �zW�_���~ӿ�
��_1�jg:s9�d!���ٷv�ʐ:��N�%ϊ5�SX�]n5=J���fa��vflw
w�G}9�������gÏX�f	�}z�O�����մ��$`|�]dP�x��� ;Tꇡ�?���>��������N�m�\jz��_l��8@��I	�r��q��;��j���4�>�y���h���o-\��?*R���/8'������?���#O���亻Լ���o
���yhQpⷼ� �����_CMGM�m|=6�y�kc<�F#h������< HJ��oۣ�W���{���� j��ZƩ,��Ow%͔R����b!�1�W�k�_���M���Ė�?��ܞ�Y_B�,��P��K2��jJ�;�<W�׈?����R���� �"��'��[	]�7C�JAa�,$������|q������ka�/
ڋM>� M�m؍�f�G�Ň��H�
=��� ������GW���A�otk[}"��P��62F�na�>Q��8�����V���[Z���bi�@���x衁#�r+/��o|o��ߋ�[=��uE,�v�0EN�'���� �FF~�Ð�)�GN���2��u�O�1,���R�즊gV�'ߩlB
�$�|Ï�ګ�<%ypWQ���d+:Dd-��)����Z���� ��z�q����ׁ���sc��' �~G�z�o�BRg���� �&���1�����'��X*��o/x''�f�����&կ-m�3��XWt7+�{�3���dp0s���ȕ~l���r<��?�2b��Ͽ����ҿB��>����A�/���qj����s�0�#tEdc�A��H=+�����)F��<)���YZ[G��� "��e�9��#�}����%��}���&�7����֭�����MIc�����\<�qV>,~�������ψ�f��-������m����p��n㴆=y�vzF�T}����	��;�_�������s����67i2���D�r��$�$W��G���=��	4��?jpKk| �\Z��)�X�Dy�� �G5�/���?�><�K�<B����v�5ƉY-�8Deܙ�Fv"������Z�i���V:���,q͹�`
*n~�ߔ7Ӛ�pO�j��h��@>h���/�ng�.��v�� �d.~\`�����E�=?�^ �/�-N�j�;%�UVA����:���/���Z���~"�\^ ��1�CP��KSnU��egq�' ��z��{�<h��x��7�|Wq�}E�17�A]����z��@���]I��-��b�5y.�Q����#�g�i��Cq,��F��2��ی���З������H��rдa�E�I"6G�q���s����o�>#�~)E�['�=��w�W��� $�v/�6�r�d�z֗BZ�tbHd��g�� �r�?�i��:�4��q��}k�.?c߆��"����w�H�ţ����F*�5�|~��4��  ���Έ)�;n⶞�k#pvە!� �ӐGJ�;
�Ǩ�B̖1��H��a��,�KR,����U8�}�Ͼh�f�ws�_i>�4x>ש_�Jicݏ*'2�� *�8 ���n���?����7�U��$�'��;�q�Z��Xʆ3+ <��=N2c�m�]�u!�k3�k09U+��i-Ηj����pUw~5�~�_-V[럏zT���y�iLІ?��t�޾i�W�=kF���x_M����:�I��}�XeE'.������#��Q]�?�4��}�<K}d��V:�R�i�\J�c�����~��k����?4}o���5���K'�b�m�{a0�cgx�#�8���$��g�U��d���j�����p*��|�K��d�H��b���u���񶿫� e͵�ky%�/�$e[hf�8ǽgR<�J����Q~�~������ �o�?7��K�{#m=�~N��	�r���V
rE{����������W�jZ�g%`�"�!��4{�Tׯ5�~;x�P��^*��K�� 1%{{�sm.���dz�ֵ5����֭w~��V�O#6-m�6��#�䪃��N ��s�@~ֿ�|O�%��/���lv��Ᏻ��+13H��L��g
�|�u��/�Zx-u��-r�q>��� �Y0s�Ǌ���ğ�T�G�Ś��������f���j��O-��Z�̹�;�uL��RH�V�� xX�>��Y�F:g�t�i��6,�P���21Uu��`瑊��7�
�e�MC���-KTV��93��Dct�C���ʞ	n+�Ƶ�dU�dS�c������_j~��<n~������Pkk�_� �I\�n8�N	�)I���c;�^��������-n��e�iIPXcԫ!�c�x��yu�Ky���^�i��I�7�f%�#���N������{�z,����}Oᕓ���˩��K�?�AT.���6z��_��:T��@�?t�Ӂ��=q��QM�]�Q]�i|7��v�4�曧�u*�h��7m7��Ȅ��*x89�\��Y����ݢZ�Z���0G���fM��|A��N�8��5���x'����g]{ŷ��f��Qo)T 2(���?�k�����0�����7����ѵ���U��Y�$�@��׭f��{�s.KX��E��msC��g�y/"Q*�9q��<rO����Y&�u�_���2j��+B��7{�	�9 �}�����۷�������+�fH�X``��Ooj�/�~2x����]7�k�dͭ�7P�7�w���\ Ē�ߚ���Xt�-O�?i�Rk-H�~�k�O>�$��r\yț#��@r2y�=+�㍕q���zu5����%��c��Os<�i�L�[m�o�çJ�� �Ś&�H�RN�O#�Ʈ2��}��y� E������}_����������>1x#Q��<7>�M{�0�B��gVVc����`0I����̰4��"�FK�ǩ��}�᷄�������5jp,�WzN�i���
�̑�V� I�4�$�Ro�� ��������+���AU��&�<{�|��Uj�V ��0|� Ɵ�'����ֺ?�/ � mjw������ń�u�pʲ4��7���6��������__�^@Syt�(-�p�|$j�6�r	���� ��v66W��q�9���K���M��3��������'�����o����n�i⩼l���G3[۴`l\ d��ޕ�~��.o�X藗I�H��l.� VO���+I��WƳ"H��$����A��:���	������^��a���M6+h%Ԃ�N��0��Wpʷ<qӽ\t	k/xV����Aw�.���2�o�3���b�ݭ�����$�^3۲H��]q����׹�D�W�KLѣ�������
D���R�Ebw	�pGC�
�ۯxw��}ցg��Z��f�.tٝ���B��rOS�U�DQ���L��S$�͝������?m��:U��l��!hf�7�x����N��jɯ!񧇴�e�u+��V�|����lx/K���^<�-�V*ݭ���n���v�J��`ܑ͊��^�w�;�~֟t�Z����N���v��!��'䮓K���N���j⛅Ԛݜ*���^���U��A�9=OC�]%��t�4[k����1���!#I��q�q(s�8��j��2oIw�h/����ͥ�/��1����I#����⇎Ss�x���+���=:�
�߇3\j�#��X+�Ǯ?Wg����l��+���*g��̱q��C�<qq3n�^�(�o���T��~.k;�%���$$~���oN��Y�������r�?�Y�+�����?�a&ՔY��S��>������_�ά�o>�0k����w9������%m S��G���`�Y��)䮥(M���_K���W�N6�L��+��`��N틷�:�Ɩ�ǬQE05�ߴΟevt�9$�X%U�2y_�Z���_������jң@�$��U`��F�D�mNBi����ݮ�Wkgü���3����k�x|amq�x�O���Eyج�#��%s��F�OǛ=R�K����}�i�u4�|�,1�g��޸�s��xO�qj����E'�%���NIS�4J)�'��3�z6���Nۦin;O����>�[�+�k�?dY�x��Q�6�={g�Z��V
aV|���_�_4_i��X	��3������r�s����L=lF.��OTy�7���ƿj�G��?���x��;ۻ�8���K8�Ǟ@�I���߶���o��RD7�L�y��Ɍ�אx� j�GH��׃-�q�&���Z�X"�gЊ�����/�]�,���6m&�p�I����ɂ8 �k�2l5g���9b�?E�vXSM6����C>.�F�u(��z�G8ǩ�U��1�i������e1Ȅ����=y��t�"���_��P�z�Y�,{|7}s=�R̀�&ѹX�=��i	K�UWW?�WN�q�=�����&ӣ�Q����0 �aY r��9��k� n[�޽E�� ������ 4Ԥգ� ��_/sHF3�Cֻ�?b�����S:����G�r�k��|��"p�[>���aq����ti'y� i�����Ht����Y�Y��j�ܞX� �t���Ǆa]Y�V�;�/�	
es�:b���w�q�?����F��
$��Xv3�@�995�2D�&���!�3���@
�8�0+��/�G%�����1k���W�x^��ؼC���z%ъ�1$F����{��^�5-7���ӵ9��n�mp6y� ��� h�z`�9�kW5g������o$�˗ ����lV� �<g�[îh?hpD�]����,3��Oá����4�{�#kS�co�xf��r>%V�E7U�a��'���мp��~�?�:Ø�#�迱�ǉ4?�ĒN���t�0�v�ߎ�����k�4_|@����彥�w������6�xX�~Z[KW��"�)}Q]�H� �_|63H�]��+[n�oHߵ�øs2]�PHAl=�����7������ ��'?�Eu���ٌ.c.2�K`n�������/Ui���ʕ��I/d�o#�?j���Ě��"����HT�'ۥ'�|Uy�-[�R,��$��g˝Ue#�=pk�~�8�4�������~�.�y�o��܎�������4��G�W�4���i:[��bI�_oDo�|�����{s�����U����?)�����T��{[�μ��.����%��`�h߿��?ę��zc��0�D�t2j&#�]}�V��y��_�=k޵��;�}�+]km�E�G��M+�FHưҩ>T�܂� ^sY�w���x�ĩ���[�+��I>W'�_#���=��<$�߽s�X74�e�<I��-���Z*�>�� I���:&qU�M��<O3�: J@��ľ"H�G$|E�G�2�u�� k�u8a���T���Z3�N��'׵5���(?y������|� p���\q��<9C�5'��xST���$x?� i�ece|Fַ��6�=8�Zn��j_	uٴ=n}=���pzI���S�<M,��i∓y+������_^��������j�[�la� c��IG�-ߠI)<u�[{����i��%��7��⨼<���p�i���=�`oت
�{�sǮk�ࣾ$�ռu�m
�Da��]A��s3� s���}+�� d��R�_	�A�j�����`m�Pv)1�V^~d<����� k��Z[�Gv�M�vr�n_0���7W~5`�>��f[Kc���ai!�X�N��&y�7�ӷ��0(P�i��>�{1�9*��{��{��������U�O���f�pi�c9;@n*�۝c\l����T�I�6*pNVq��M�ʒp@Z���w��Fx8�R�lf`�D�F��@-�ٔ�|��v��)�iP����zm� U�pŚ5Ys�åE#yr>T�Ꮤ~t$K�#;�:s�YxdhXĩ�zn'�֨%�W��|��؃֮&�m�^N������x�D�҉ �$g���G�׊��v��X����⽯^��0���H��܃n`U#=�g�x��s�̩F�0�4��~$jO��.�=�kMa�Ѷ��+�3��|n��/�(�Wٿ4����%Wñf�η����n��䐟��|e�� m�����9�J�#��&�O�:t�_g`��PTJ��6��q�i�æqM(�8��{O� <�{�\S���'�L ;S�
���w`ƌ�R�ޚ��( ���@$���
9^�)��ނ�6���Q�<���4 �q��?�+�

���{�N:P+`t�ړ����q�8=[���ǌ����~��)`G%FJ�q���AH���6�5��?����3j����r :���\ �S �׌~�����~��~���y�/uo�[#�z[���G�dh��I�q_H|����?�c\�M���������X��B3�q^e�E���O�H|M�x��o�O4w2��4>Ғ�f��W�9n9�OSX����_�� ٿJ�w�+O�M6��z������<�G���n\��|��������SB��N���V�E� ��X�4�B5��un��[Iv�99_i#�5�?��ſ|w��4�Uu�����AH��l�̌n1�N;W�~.�=����i������^�����R�]!�p�/�w�Oj���M��g��UMSN����U��I�:,��~@�ѕ:���z
�� ��?b�3jq����$�#���[.ҹ���|�3� w�x�*xM#����ȉ�U��g�%�z�� ���N��?�wƞ�]�4�y�E�Ey �DM���J�F\���s��%���?�w�.��o�Ь�����a��̳["����
$,
��@�|���í}��Q�ԯの#	rг��M$nd�!�`��(G�?H|Q�j�W�⑱�^�+x��"����rY˕�J��n�py"�.�_�R|A����mWU��O��Z�������!yрX'��V4�{�Sݵ���%�,�:��me�36�7��;�
�����%�)���v�����j��?�W��}�ۭ�����.��<N��!R�7��9ϵ{�����E��[I�W���G�����7��`�Ba��`�z�1ּo���ƥ����'�<M��-s]��!��{֙�F�&*7�Ĩ��{	�ӻ4��VG�g�<i�oi������i�̨��+�v���0���_�'��m|G�|_��/�,��DQ�l�G����== ����Kt`Af^9������9� �W�[x��w����=R��Z�UYJc�xs�d�%78��[7es_C����Y�������,d��4qyc�پmc `�r�Ҽ���(�j��:�Z�ۼ��*<A%HRc	$���` O�׾�(���.�����4������o;0f��n~�W��� h_���<�x���ӵ���._�>Y1���-�`�g>��-,}��L��_���Ig��XS_��"�$0�%�w�����C)PA++�g��<{� ��f���Yﯖ�F﹕M�eU�:�q�`{���B�[�ց��}�x�=me1���S���|�Cʲ:�ǎzb���� ����9w�gÚ����Nhc��n"�S=ҹ$q��#9�Q���I_C���Bۂ�30�SF̫���k���������{����O��c�T'd�p�;�~����g�?�w�ƆW�	bf
:�߭�G���i���Et��o�^}�^=��C���|��m2�Ộ��~�$*�~g�Zr���B�զ���!�T�̈́\����=k�O���Y�_�wKҼu��Z3�^xI�d۸!R] �p
��SԿf� ���y�V����o�y��FO@�l��j����?�� �(<i�闞�M���n�F2&p�̍_ti��F3��Vr�jȸ�E��?¾����LM�5��m�N�Ds�9���I����q�������}g���c�_��Gh��;����r �}_���?�'³se�X��D�������Oi0*
��|�A$�o~���|L��>"�k��N�v��I���i���2x�I�>o��^��)��ί6����o�|m��w���cػ��D�|��>A��f��ڣþ1����ӥ[[��e��6���/`�Knt��ͤ�n��^KΈ�����x�J������;�//#�"���Y�yyl��I�m�/�O�'�[��R�|?��֩�( ��]�� nϹ�gԥ��mc'�o�/��]�S×~�+�{�˔�@�� �%�8�k�#�G�|P�>��C�Z��;Kt���XI�&RKs�����m��|O�Mz�K�J�ӼD�)���Ir�.ݧ��G'>��������S�4oiZ��/�]��~�u ?}�j��F@�2N��&�EOM�� �
����~��L[�=
��V�Gn/!��iJ�?xdg�|a,�Lb@�sq!	�]�� �>�Ҿ��7���G�b�Ń������	t"��oI摅�8�o�>���S���(x�A�� 8~A�=�9��T�ʵ���x'E��|>�;��ng�u�	<5�d�1Βm�Sm^O �T�+���������j�w����s\i��G�f�ޠ�1��m�x�H�C��<TuVK�F�i����r�U���,O|d��9�6xv� N����0^Z�mu����;�^"��Ͱ�}ݹ'�je~�K=CB���a���\�����[��̓��wU^�<��Fާ5��$�����BYݘ��r}�Y]�Y��F��o0�#f'��������_����6qL��Rp:w*F# ��ҕ���@1�^��<���\A�C$1�$t=�N�sU��#`���� �⭸ w?�q�L�ap܏�)�[���l�s־��M4K}y�����ubs�׃�#	��?�{���Ꚛ� �cÌ�i;�5�� )u	RO�����k�ʑ����sM��欗��ZA*�6[)Db;��kʵ&� ����z^?^��)K����דQ8�ٟ�b$���їPA�,Q��8�*��<�kt �Y�J���2���^��­����=O��'9]�v��%rJ���9�\b��z�����n���:�c%�����6Gl�U�]6�Gx���ƥ�*��g��W��˯�	�� �㯦��|����r�gS�� ���Kҽ��(��(� q�>�(���(��|��Y�oZ�.��ã��&�i��2H#�oz�|W�~К%�b�$W�e���[y�d�B	{��T�]U��c�ύt�#_�<H�����>yX�����C�8�O5�?��tA�hʋչ-</���S��&�u�'V�Lzn�%�2*G��[��NH+�}s�׊��Zmkⶽ�Hۖ�|���a��D���s��
���ݳ���|����Glf��t���Ip����>���_�.�YH\�{c�澉������>&����n7yS�2 E��=;�_9�f�,��$�{S��4�:qv���W�|K����HZ��_�t�l@�/�����)�4�դ}��N%��*G�+��|L��$�`k���p���O����W�� �ǀl<;�i^*ҡ�	����EM�� Hq�Sӧj��>�>���K�}�m�OC�S���jHO�Y��z��_T�F����d#�>MǍ��*Hn�P�ln��GlI�_�#>�oq����i�+S�8��o�>-x���Εckͤ�o����6ye��?*��O�ī�E��i�X��,q�l����>���G��4�5(�#��3����1�_�Z�,���n�|^����[춫�?�n��ç�S(��"�b)�z�}�]��~����c����s]�O���L�i
�˓�iSvr��=1^��/j�;���=��0Gu|�>b�$	��R{�T�[��:c|P�k/lw�
�ݜ��}3S�7����o�����O�ɤbc�O-Q�� �#��ߕ��:.�Y��U�f�N�5]X�ه���[�^h18u�V�˂q�XU]�S������[��֍t� �V_*IA��w`���L����� 
�'m�U��_�=�%��-� h�+tb�/z�y�� ��w��QR�od֝�y�Tc)+i��
|!׾�yy��h��a�J�d*�y
O<���~����2�)��d��ՙ��`�2G��� 	�$���mu�]f&�g�<�pq��=�q�f�4/˪����pgw��kp�d	ϽrV�������Xl]/g�h�۩�/��?4.��^X.����U��~%���e�N��.v��k��Y����n�I��SL��\%͂<RH��J�=��k�mu�y8l��W��+����E~/7���p�U�����W���x�>�;_E2]���	褞�Z�j_��α�~MgJ��/P��Dֱ3��B��#����ߋ[n<M��~s;���^��0����,��Y@6B��'��n�I��~��N�RI�cÎ*3�u�{��φ���2x����w��-�-c���TM�F� �}*_��:�ϊ|�_�B���Zn�%��R��H���%��;�h�5m_@՗U�5;�MI?k���bI�.H�N=�{�� �o��,��_jd�mZ@��wڠ�s^��\���V�_�KW��H��Wð�Y�����ϣO�r�ʦ��{�9�����H��kE1��Y��|f��I�;=j[�NmJ$_.� C2�8���k�����X���d�	%��[�"�T��$�ӊ�ꔽ�ھ����%f:O�G��C�&��b9��>4y�0�uٓ����xg�z����#�Ě|>l�Hg�!�T�|v�kR+����7>[]���]���*!*�:�_j�k#I�wr��i�?y�ߵc*n�RU4�{��SP��x���Uu]Ky�i��M�b�r�o��_1�d���,x���U�k���F�+��:��8�TW���G��-�h�����ӯ"�F��Ӑ���(/���.����I��-��� gj��ŀ�<��'�(�6���ѧh){�W��l�ǆil�D������R5�y�ٷD�J�ʰ|7�-�	0�z��)S�����WM?�J��s��>�jf�@6��v� 
��\���,��5�qoef�G�����5�,�Eȹ��z���έ����U��=p).-�$nu'�p1[n,�=��s�FsӷZI�D��`#9�T��@6��r���8]��=�nk�L� ��V�~4Cf��
�m�m�j�Ê�6'�c�����e�]�c8e���_J��\�L��e�ڱ��A�i���]8���ʁH��Y�h���*z��� =k��A����9n���u���>_&b�$��2�|�i�7��I�6�3gs㎟�R� �'��W3�*|��MMrA �7���|mj6�j���}�쯈��P� �.~@-�E��܁�Cy�6Iǰ�_���!��`J�p=��^������愇��x��mf�5ڢ����pu �c�O�#_��X	UH0,�1�}�oc2T!y�C�p2*����1� #$�Ӝ�ޞ���A����@�w�>��g��'�x�]���}��c=��b�j6�)�T��Nx�G��:�K��U+ч'�@/`. !��s���
�;�1)%�e�� �9'<p)�1����ޞцR_*L
�u$���3�H8�}��L�hk�Y�\� ��:��y�JC%V�00�Ҕ��勂O���2�IAFR�<����4d�ρ�FF9=?��N�D�XG��k/��t88n���!��>ly$߿��-�+�ެry��^޴�{����|E�hWV�Y�w�Cnr����P��FAǯ�zƽ��W�d���,%�r-���Y��	R�+�k8*��� Ǌ��!ǘ�<WG��↹���o�<1�ɧ�2���&�<2�pU�GL>{iajsڝ���/5���X�A*yHz	3��&��0�E�m�$�n�$	`mFf$�A~ߝ{���p��Z���S������[���4�Y7�"�E�^�*��\���=�ƞD04nL����X�2'���~�R��ԧ&�ǐ%fy�i�||�LY���G��Q�l]D��K|� �N'����^��9�yvB�8�H���1�����x=�͑ҙu�L]�k$b�RyI�IT(�!<6�6��� �MF+�<ϱ���oQ&�9R��s�G�<c��9��Hb�
�?x��{c��G\q�q�׳?�+5֓�����v�ב��Np6��/��� �ol�-�Q�x�r�ax�;��U������
9#t�y5�>q�b��^XC����s�\��,�9�O2��w8��q�J���_���|e��LOɧ�lV��^7��v��C!��g�� �G�����-?TA[�bRT|��p�G5�.��7�?>�P�{PM��y!���$��a�XY�\Z3�[]Ìe�q_��� ���-��!�����k��.#�[c��	 �����k��#�Ŏ��?��b;���Kb�������q��{��%�R����%��I��(����`ls���*	�co-��6ǹ�s����ϮE~���O�	�d��Đ�8�`����RP�F��vNzW;�C�
Q���G�l��C���g-���`[y�U�e��-ܑǽ	ߠ�Z?;E���I�(�B*�M�� ��}��&�U��.&O(��ʲ�+�>c�Oa�+�K�?�Q� ��"�݆�íj?��-�ye��
I`�N��t�|�#�O�����iuwò��.��6��6\��W����$���Z�������.$hfydf��GϵOq&���0��]�.bc2�L���y�g |������� �Q�\�M��-��\�Q&��¼r[v��'�����kO3ZYZ귞8����W�`X-�@)� ��T99q��rvbvJ�s�	5MA�4�34��os� �@9�S�&a�r�q�xO�M{�����z��i�$x�d�b����ٍ˟m��zd��6�XGc`�L�GS�[	VN���=�WD�Ԟg؟�0���'�Y��N֬WY�n5=�Ԅ�`�Q�N8#8�=d.�)�=��-g�Mψ�5�`��焞Д�|����w�:��_���π�a��:E��wB��)4�xٟhRDU��a����C��<G��k�~$�h�<�������n��0>h�7�z�r��������������r�Om��V����kMb!�]��E�Q1Q����L�s��P8!���ٕu}<����Z�۫6�-,L�s��<��^q���*/��n�u��0���K�x����bX�@i���=k����{k?�i���X�׆n�ҤY4�n,͢�RQ��	�{����h�?So>&x�� ���x�H��$��2x-�Ai՗#���A^����N�|*��>�*	�A���Xm�d)m=����d�<E�?o+�s�v��1�)�����f�;��ˏ8�� �'�5��o�
��"x�g�]�\>�{5�ܖӘ�e�	?�|�.w qUgk�Eث� ����1�u�xu-KB�`������fX��9 u>޹���<j^���:��[��|;�O�l�ƛ�iтln�T��c� ����8�|�_�շ�5{�9�� 	i�A�;i v�![b��0@;�C0�z��j����x�~�u-?]X�O1Lq�S��RQ�g��!j}��0|r���N{ߍ���_�� 	�4�K}
��ݜ|��r_��.Iʀ �:~?�D����Cx�]���kZ�.�`��d ����F�8�'��u��*_��K�[�Z��]?T�-��Zm���l����4Ep8�xſ�q�M7�^0Ӵ_���&��]5֙�i�[K�F(��LSV�w��a�(��eե���T�ob�.!� p��:�F���� ���>i./.乞��g�c$�3;�z��_���,���R]\J�M#��m�ē�I,I ��$�{`P��c�3m���r��$``����R�<��'�}�B�I9{�_5v���z���ӥ*J�W�������OGf+)fR �S�#�n�X(�;G��i�d{X��m�>��#��S���>��af�x�sLY"fQ�nf���<J�F��f|������$�K9a��Q���׽|)���]H�T3AMxO�+9f�B���F�� �]��L�"� ��?�L�l� Jqg=�÷�S.F>؃��:�&[���:��y��>&0 ��==�zN�,�'�=��^eW��#�lT���YG�l����Q�H#h�Ҝ��/��6�y��0�rwOҧ��򒽐�%P�v C`縭��P �6a�}*�
>Fa�3Z����G��Y����ҽ�Ϲ� `c��S� �J_�}4����G��~L�������^��^�t�?u�� ܩ���*�h(���P^K�EIj|%���[�I�[�4�_���}z���J�G��֣��Ų��;�o-牃2�W���KEsգB�8���k��DУ7��խ����b�'��>��⚓jz>�����2�X�������2�T��b��_Gy�i�FD`r1�r9ϭ_�� ���"��oc����D�H�dCj��	<����������x�iRz�&qږ&yx]�`�S��Wҿ���c�φw�{�o�ۂ�ǿ��9�zW�_!����C����4�]/Y�o�^2y��c�1�9�zW��XfTy\��Ǘ��3�q����������,�#�neVI�
�sϸ���-�G�xg�:;�ަ�!��3���ڪއ9?��y��ů�ڥ�Y�Z�(1�0�8��\��5ï���h~#��Op���';��7|z~��9nKS��|d�g��Y�R��Ti��R��#���i~�T�uxT_���������5��_|�x�+xu渶�NV�g�\���v#� Ǩ5柴��X�T�d6�\ǩ�ڬ�޳+t	���������/�mM?U�.�K�R� ������1Ҿ�6��yz�
�/n�h�� df��O����*�c�Q&1��Ҹ�����>92¦Ut���˶~���ɗ��<M�K	�F=ӷN�����l$��a�f� �1��J���\�l����9ք{\��-�: X�##�|��lXķ�o�&9q���?ʾ�k��b�1�N����mfj𢓒^��;�d匆����ܾ�K����ƚm�ّ�!>¹W��� �ͥ�0�������ŏ�}���� �\�ę�å�$�[�~"�J�w��E��N_9��S�Ѵ}׬X���� Urp@���H�V?�~'%p~�3 �`��uw��]H2d�On��'�3�� �[‑m̈́��?���)}f7��S�J�;Е�J(��i[�FӞM�� �]�ؾt	�j��Om�FA8^O��_rZƟ�����<0�� �ƾ#�Ζu�R����i�w��D�ݹ�~ߋ���'��z�iK�S�8߈ZN��x�'����ll��paD�Iv���K� �2L~&'��F���_�/�jg�σ�}WV+j�G ��6��}k�~3|=��_�>&����=.��r:U�+ǭD��Լ��ӣ��xd<�s��t�>)�o� �y�O�0y��<� �C�	��"�y���(�,��;�d����J�����j�]4�ú����V�5�ͽyw>j0z]�67�:%φ��a�u8�V�ƒ6ɣ�ˆ}3��˪7�'������\���<��4������L�]q��M�ş"I"a��<����t}�G�����G���}>�l�m$m�-��[��J�٫u=qi���ڕ��+�Z�B��,��sU���֋��`��ҥӒ�&ݝ���sZ�����"kH�מ�3�wG���m�<u5_QӦ�滺��IVa�VУm�N��^-��U5��+�ʟTy���ψ5�왧�N��wH(Ɍn� 
�յ�����ɒ8g���%\5��k�q؜d����>�[�,�j'��t�t�v�y�or#`��s�5|V��ύ��Y�5���R%����*��q�{|ۏ��a�
�I��O�xZ�/�g���k'x���ݕ�roo��>���ۈۓ�}3[����|]���>���6x��U|������z�\H�:LYy���׳��?K���h����m��I*���*Y���H��xUc���7ĞN�<�}�n��jߵ�4BB
݆�UfY�O
B��Z�9#���A ���C��F�6g;�������GG����p s�I�2�h��u�9=�Y�T1���ן�J��J�8bM�ˏ��:�I�6�|�������0;IV4�0GӞj�w��Nu$E�"���,v�,A�9�����G�خ�ܖ��l)�=�v��g�#���+us�6�p�=�¼�K���ǉ���;ey�%UH!��q�1��\���o�L#�̷�R-�/�>���υ� ����-�O/�n5� x���/��B��Y�X�@�r����T�I#��h���͇���~���V�bԭ���"��8H琕yN3����\'�>#�9Y�ѵo���SPy�V��p6��e�+n�<� Ҽ�A���+ay���*^�Y���c#�[��N�9��䵖�X���=����Ts�2/�1?�0q�W���s&|[α2��鿢�|/𱵴��&�9�Z�aZ��^r�&A�>���9���.�]��~�)~h�ܭ��S�n8>KHwG��ʞ1����,�O>�M��iO�|�g׺�ݪ[�n%��"�c�����ӣ��z>?�g�ʍ�cE��}OV����;��=�����/�d#\c!l��0�{��?>[�V�O��;�]@n�K{y4t�(W�ar̀�~l�� �_b�g���7�؁���?� ��� 
�5�9nA�E�ۋ�M�1�'��� {��KV�Pͫ�����J�E��� ��쬳�J�L"6�ځ��r �U5O|7�ƭ���?�~�P۞��#�c`����N̤^B����њ�[fߞ����N9_J|�.��=U5ms�R�,!�8���zcӎ&���\sJ�[���/ x��n�>	�2=�T�mc��D�5*I���>�Ms:���9.�;��:]�m�-�B���8��m�;㓟??t�!�oF�`�aۑۥI��>�N����}U�F�p��FX��q�Z�V��Ʋ��ms��G��j9���]0jZ��$�.Sc@g���v�x��}������V1*jH�M%�������X���I�W���,,�6���ug��3�*�#j�>�j�l�/dxUᮛ��i�n��1�ү���� ��������i�m�K��"����fR9#=)ɥ���Ťw�5i5K֑mjβ��v�(�H~{��甹wI�/�0�7˥i��\�}{v�֚=��Ա�|��λ�=H�����Pݏ^�C��� �Ԯ��t�W�� $-f��1wj��ލ]������ۯ<U��g�������!��u�V�ui�d�8=��)-!ӠH�/�E?�[6˩ˀ��j�Z�w�[�D���;�R�	��-�o�wD|)�}2��V����!�tW��{�[���<�t�|5�:��\��'�c��_���x~�S����5�-��ԥ�~/x�Lc�a��Xi�i��3kv������^c��9�8y�=n��z��_|�m�B�Q���9�5�:է+9<Ҳ^����ψ�t��$Ԯd��Zι:@��lO5xm��#��]%Ɲ�7B�����R����k��[˓�����H�zdc���W?�4�N�"��u�>R�tR�Ӻ���{��Yqi�x������>0�`��ł��d��͕���]���Rql��8�_����M�G$qH>�)d`�u����� `H�ǽ4x{�\�.?�W��{(�)�}ۉ���ǧ���Awf�\���U���\[M(��Ht<^zc��}b��뿃���&����[�E���2��r)<����a�NA�jş�� ��o��n��/5̆k�q� ��>e=jΥ�K$q�r���_N��3x|�t�e@��#�:qN1���� �If���\��ߖJ���">8��=�ךև�� �-m�<�� ����k���Y����9�f�YK��m�<m)�t ���Fi����}�����G�Ⓧ����?�}:�������hLkouq3,��T��.;�^9��n~i���N��m���V�Y
����q�\��񟘬��8�}��;I4��72�`{t���ٔt�^|Ķ� t�)��+LXc�g��0H+��V�"�Cw�Cqi���Oo�<qy�S�q���s��Lz\в�XJ�*�G��O����갏��Q�}3��I�&�?�MɧAb���U��۴���v��6�� 8\��.��,�M� 
��$�#���'k��a�d��n�FI�e6�����e!����:T��I�7`c��9fPĎ��T�y�oK� ����K�&��U�dg���R� �:aO���r|U������M�f��jP<e��{OҎX:�$3s����8�,��D��/&7�J �u���x޿���3��������0=��V?���3�� ����!��fi!����ܸ������o��t��4)m�fΣ�Q�!�`�I���H���Q��cF�lL��2�ը���;A	ԮI�׿��o~�:���kk��S��٠�Q�d�"� �����.c��E������k���v��մ����1����^�`q�N:��������=��E����1���I\��
�=Wp���?�>0�|I�6�� �&hV>!}.�q#[����H	�"�ݖ�ry�~���>;�σ�ŵ��~�r�1�sF�������Pk)^�ѯ9E4r��?]�-u�>���D+�\�'��x����z�^q�πP�������� �Tw����lÎCv�^�g�W�+�.$��_ 5-j8\wn�S���N1�W����_��"j�����xgGgc�fӣ�m� Vx#��=�:�*���׶��m�t��h�Is���դ��7������M��7C$���q%�Ѽq�_̶b�V����ϵw~����i:v��ٺmĊ��o���d���z q�p+�����28e���5��[�M�-�ڶ�6	�<�U;]ȟi�ݳ��|'�'�dV2E�m��DXs�v�:��'Һ��W�/^ip���,Ҩ��P2ȑ���9L�����x��_�_j>��A��Gh�KM�!� �9�>¾����^:֣�췶sY^�-�YJ�E�$`6�9�ϵs���LFcV�Mj�u�?c?i�?��ş�����V7Z��bE?��`���8;��~þ��:�7z��Z�P���j?�;�Dʥ~nT���|�^x�Z�o�{�~������<���6�z��'��w��}��8�MB�/���k4�}�ᐩ�`0�N(�yӏs�~��x��Y�m�߄�>)��|Cᵷ�T��+ݷ��9Q�'O�'�~�����{��>��^��~3��5���)T$�0Ã�A�?�2x�mPI�=[T�� S&�4���c������#�����K�+<vGV�ً����!���+ZU}�����u9Z9[��ट4���5�<�a)����I��X�¶�zb�����?�!�KM߼hd-u�����yd}�~;�?�'��(#:w�kE�e�&h��VE�8/��{��+/�GIo4x��^����)N���=���C�d������s�'�zQ�N��nx���?��?�|M`�1o�W�2�\�cm<��6:�+�� �O�/�:��������6Id'��XZ�PT��oB�9S�z����������x�W��4�@���i��AfVV��l)���$�� |���?���⯀��C���~����Mzk���ud|ߌ�X���4j����+��ٞa�x�g���<#���[^�Vk�{��p�_��H\�c�ɮ���7�6��B��dZv�����y#���j��WR��plc�z���jW��l<m���R���t���>�iZc!>ᇾk���� d{���ŗ:��%��4;11V�͖rN?�4�匪�*V>�?��>׵MS�|B�ƕs-��h�cvV8p� ��;u�?��uM]bg�%�I 
̠�	���|z���Y���z�σꭨj�9"$��k�&�;�	�c�W�*Sz#��aU���� J_�+�5(J�N��pz�{~&���S�
��� H`N5�T�`ϓ�K�3%a;F8���2˦s�OQ�>�*���"|H�������Kuxڅܷ3��� ���t<vU���/�]tf�/�0|�?>*ۼ0����2���$ c�g�����zl�����)�IΣ1� �R��^��_8~��n@����:���5�tG��?��?A�QEQ�5��֠�j��҄^x��v�B&�r�b�ˀE}vFq_&~�.��_�f2~��Î|�i˲81�S�RZ]Z|�6�o���}�nb�^Z��>�?P�7���^���1#��[�����=�[��RY{z}k�o|=co��#�S��rqԞ��.�a�a�օn^K�M&�����|a�Nx�>�>��G�O=�$��r��|��mf��ҁ?v�^��g��J�9�n�����^��H���d��\�.�����qU*t1MR��[���b�����f�H��(��qޢ�s�q�Ƭ*��� k��[�&��h�g�6>�V"�1���D��?�3W�J��� �eቯ�NՂMy/�=İ$�;�{�qӏj��w���2:TW�l��.��B��cQ�J�cG���8Nǹ~�:��� �ږ��Kv�k#<IC�v��9���A�7�x�-v��au3*Gd����9#���t�
�$�|2׎�ii������@=I�J��� �wM�F��RI�W繊N�督#��j�R��º�k�C�|d�Þ��?m/����r�p�b�� ���h��>����>����~����Y�^����:��:o�|
����9'�H�K�+���^�Q�pG��U8����/�`��#R�w�=�fi[EШ�g���P��bK <�?3����<Ee��K��g9���)N�2�q��<W���UK�� 
� Ep��I?�!p*���QG-σ4
����G5�*4d��~�c��Jtk{HKX�3����+H%]'[������o����#�^��G�k��uk$1;B���3��]�~�BH���\�R��8�T�NqTn?k]#������H�>�A���ѩ�3����>�R
2{�ܡ���&Ao�K�T� �=|/oUA�d ��s^��ڛ�8Ѥ��]/O�����;YV����p�۵x�q��!�;���ױ������Q?8ϱP�8Et%��q�|7�|T58ws���"��o�>��}}��5�����/�NBGOO¹�����^8>G?��v�1� 
�E#j�;iT��sƕYԧi3�*���t���hl>�)�T38F��x�`�V�-g�z֫�Z���%�&��-����8�K���\W�<���K�����ߵ$����s� �G'��Fi,l�O�}���ܲ�:�rc��zs�M�m�(�t�t:��{�V�!�K_O�}]	��ym�P6��Z����%���k�U�S�QG�q>[�o~��NO����}���v>*DUW�g��� zq�j�����M����O�B� ��$ϤLy��#$�g��*.G����WhW 6@ɿ�� �Ymg�Y�6��W1j)���� gڞ���۫���O����KO���J��#���5�2���%�78j�:6������w8��,w*�ڸ���6��.+�y��<0�{Th�.N2�.��=�գj�<�@�����c�H����J�4:�с���iI��=1�t=������o���{�#Ʌ�=sUsk��X��/�ҴQv4w�=B�uM�w��>�I�S���EW�/��i�v��Ǟ�����~:|�w���+�7[�it����
���Χ��5�L�Au�����;���G`}z����?-�EO���@���}�c6������B�3�]��צkա��Q��yvk(Z�c�km,�_[���V������H��k��߰��ͯ~�^)�֡R�s�B�V��u��8�8'��ƞ�W��r�I�^�y��@J���d�$`�G�FjKC�c(�ދ;�PZhxK�� X���W�(֎�p7�0*+ʗV�i%�:��X]I6 p?ʨ����TR�����Trx�ɍV9��9�r>��M��y��{����.5Č��H��}}��S�����^(y��vE^������j�imKq!��9'!Tw�>ս�_��3���%��4i��&K�so
�y
�u�y����7�����Zjwv�~%������a'<A�2� ���8�e%�Jغ8uy��?��	|�|_��N��E��6K5����t��O�����[����|[��/�C�k��ުt�K|va��b�**�8� �S������[�s��W��mF�L�y%�b$�������tZ�z��w�3[� �5���K��8F�a鷸漟�Օ�ˡ��m��T����i�i~]R��d�o5�m.$ �nAޣ�rG>�r��M���L�6�k?�s!��R���c��q�V<5��mt,���8�A"�Y@��P�Ѓ�L #,���$z��^UF����U�ԄmG��'�8�������H����T�G�����L��Ӵ�Ԝe���㨭�ۢ��An�_Z��e�;�T� �K-CƗ�9K�{[h���(� �����De�G�Ų��k���%� �����v)� <b���zʵ���,�[�k'mDThl\���ď2Rz��گx��[m#A�-����W�£�d|�-��������|+>�s��yl;��
I^	����`�9�4x�Ud�kCӒ�_λe�uHX�(�
3�^p;�>�g.����Y~�T��M���y� o����o����±���n�}	{X�.�f1���9g=�y�������<h1_M��n��O�n��z :(��|ֳ�*^d��96�m5��4H|�-B�B�iA�rZB[������'�X�-ǎ���	25��Y�Q�9�ֺ]�����;º��f�c�]�..�`�y �Ìp*�-�3��3O��ce�˷t6��� #m���0�n���x��]�[��'�K=KAh%�]?��3�C�� I���������^xvx��u��44�?��x}��$eG?�tR$��Yj�z�v�.��� $>�� 皸l&��Id�ֹ$lڎ�͕Ӣ�y�6I�d�^}Ώl�nq����.��ϩ�?�Z�����c�߯OZ���:-����A�fo*��w�Y�!��;rGcҺy�ln�Xg�տ���}��a��S��aԨoQ�54˩k�6~j\������}*Nm�d�����>���f��/u�B+;W����@���5���$���9��3ٷÿiZlׇVi|	�F��^\*��wg� �`��lsԐ1�=;Gд���.�5����"����ψ'$b4�'��G��~n��:�Eώu�}<)imf+KH��o��s��=�{ Li��V��&4cyn`|F�H���u(���4�u�O��l��+����9q�8�_�t�E����� jO}pPV� �#;��C�עi��K���h�^I}m�K�!�#�#r1< A��Qh�>����ǚ����#g����zWK�n��ʴ�8���k��z�wb��M�`�b��}�yv�����|)g��lf�c�4��f^%db'��#i���-~xz���:���s-$���	�?�8�^
���-u]/�_����c��>Vs��z��t��g���y��uۍ�}>��]۹�hd+����b�C�<�P���^��H�.�h_�?�?�z7�5葢��d���3�B��=q�-|��2��x�_n1�j��QM&���QU��[3��G��v)�޼�֬]Z��.9a '�q�^q���I
#8(91/ � �뤴� `�4�eF8��h]�t[��s
$ �̾ac��J�t��m� uwv8��}i˪E,1�yØ�Ʈ7�ʧ����;��i2%�T�~0v9V���i��R5W`p�ך��/
<�0l��u���X������=w� Iim$��hn{��Trڃ"�H�o�y� �R�נ�������n�����1��� �g�Y�P��x�}ߥfk����	���[*�(���Y3k�����);��W�OD�AU��ɠ[�z񺕑���N=�ٿb/�Z���O�,�������V˲�1�>�����߈z�-���Z�!�I��+����]/�'���?i��#�#���tֲi�^G%Fބc�.���?{e���(Y�ģ�# �����P���GQ��<!�~�����^�_���a���n����߶���S���W��,������^�(<C�Rs��_Z���xV���Y�G�Y�1?g�Q��!�����w��ϕͳџ$^��>������$�׆��9���:\w$ ��C�=��W���_�/���u?$z-������Ȅ��V`Ir���:�k��j�� ���=?��H$e������a�5�xW���ރ�5i���J-M�{k��������B�w� q����F1}S��p���мA�H�#�?���-a��Ov�a���є�\�����xf��cE��D:��k�xnmE/�֤H��8���ڬ�?.󜎕/�<uw�O÷~��?�c�z{���~����m�I�'p95���جP���i���F�z�F�Ò�v��p@��ZF�a�=�0�\ͣ�<�G�[�FiGE�����������w��� ��BG��|T�k򶇨[��d��dTxc�����*��kþ�xӼ�O�?�7��xm��qx����m��p��5���Ğ&����o�� ��������Z[���X�22N8���r�OA�����j/?ko��h#�H{q�62�ʜ���z�Zƭ�?ڊ	��ְ7>"{[�U�;�)�ޕ�����B���o�xwN��,HQ��`ۑ\��K=OZ�/�>��W�1m-�ە��^�Y%�$q�K����O*�~���j������B���������-4o�@��� ����5���l����:W	��/�>x��V����-�}}nt��6�;�s�_:�a=�k��_����?��Y��<q�JM��F`;`px�>���߃^�������D��v�z�z�ՠ��+�rT�2��M�u_�r�KC����럳]��/���5�ⶆ���!啂����V������,|h��$����r?f8͜���C�t��>x�ƿ�q�5�k}@�&b��� ��z���sX���G��wy�Kg�*�Tα�]C����펵��U/��To������G�/��L�n#����K#��`'RٍKm��O��s?�`f��5��SF}.�����cx�ո�a�p}���?W����]}��?���5���
�-��~[p^pA�\g���#��8�F���w��m�}>��!�4(��n	�rI�+nf�>����>2ѿd5+�!���!��Z���o��e8N ��ҽ�/�šj</g�;�]oC֬'�-R6W�X�%2@���`q��Zn����:����.k)-n4di.e�Mn%�`���O��s���/��|a�^��M+H�t�:m(jV��*p	g(�9����r���gmO�I��޽��iV�_XCtC����Xc��ʮ9�=�����ͷ��lƟ�w���cԳ$r�hd���p"�~,~���+�'�QiW���ƽ�b�>��wc܃]�G����I�������g�Kv��#�O��w�7:w\������H� h�h�
5���?�ԟ	V).�-�h�P3��f9���U� �ܷ���r�9�z�C�~=چ� Tg�s\X���\� �*&s�����t��W�_mY���p> ��Ķ���<
�;����^k����=wr�F������}*f��Z�T��O5�Cͽ�����d�L���@ G�X��cU!�aߚ���o��v�����ꎚ[y~ê��Z�sn�Ԥq�:q_C��|��J_��s���?־�?y�?�i���*�`)�N��Z ;��C��Q� 	��݈EO5�1 �9ɯ��W�߷%�#�Ӓ@&x��k�R����v:Ny�C�ԼQ�[��_iцy��~5-��/]Y���i��(�]oSq�ȯ����m~=+L�i��2��&N3԰=�����x<=:��g�Ζۣv*3�C`t<f�<�Մf�V�e���U�B<�����u-'T����Y�]�ܶ�����85�j��#�W͜�_BE%�#w�X����Z]lWٲ7ʜ��X���R����G�Rڮ�y'�׷����PXx�����U���f$ȱ�	���V��$������0ȯN�9oc��c�7���P��#�;;I�2y��܃�J��=��O��Q���<����m�G,m����8����p�[Y�U;;x9�޽W�� �]��j�6D�m&��-�[X�Xٿ�H������-񗏬��f�[�:�"V���!���0;c���q9ϵh������	�\����"��������*nÂ�����|��|U�-Y���7�=��<��n-��?��t�<� �g���a:{ig��1�������W�~�p��V��p&E>��ǘի��Jteml}�Ѓ���]@�K�^/�5��#]���0nz�ϭy�_��,����i�g�.��̋�yd=8z���;Q���_1~ܑ�z��Iɷ�v�`����yNi����:��>�<���a]J1�Ge�]�$��I��l��l�E����\�~ؾ:�>'Y�i����d�;Z�:�!rr��>�+�������?r��8�߄>����3N�K�au�´cr�Fw`�1���_gSR�7�O�2�UJ��So�z�_��_ZH��G�����١����~5�㟊>,����T�u���E�X0'�c!�U�zѭ��|��s_�����'�96��3a���s���(����IOݾ�H�V��nt��;����,�,�Ьcդ��KAdBP6���������{(������<Y����c����!n�B��E��R�ʤ���$���)B.ڴ~İ�
�p8ό^қ 	c��+����|(�G�~S�x�5b������V�w�V_�z��Ml�w�nC�>���f|H�[��r��]�'�r�=L`�=H��������.f�w�w�.��kMCZ}�O��T(JΧ�px9+��o�4Z��IФ�c�,7���KpH�u?�r���iGR�/�᝞#����X�r3� f�4_^i���U���jZt���j�\l] �x� q۞��Iӓ�ќ�u=֑����ǉ,�'��|��j�lt�0s�l��u�Y�^"��%ĳ�=,�L��� G�F�R!�
�s�g�Go�;E��_����mŽ����
�ud�v\��'k}3��_E)��Rx|�'9� ��z��R7��S�l��6������iI&�BC����� <fﰞ3�� �����������f���OK�Va��Ż����k�F��.�v:f�n<�WN��Ek��{�3�=A�b�M/�"�h��
6�1(���;sY+-���˷m{α���]q�:�'�?4o�,Ҽae�Mv�]Tmi��n[p���oˌ�y�i��t�0S��Z��v��$ׯ�T6�����C��X���Bړ� � x�=zZڄ�N�籄�jF\�n���F�G�}7Y����}|�TV�:M����R�?.�~l��J�?��i�(O^�AՓ��b���=�D�}��>z�9��XϨ~�z-����u(�6��Ȧ_,�d~vG��Nk~�<�s��Ϯ�� 	���e�E��1[E9\.ZL�+�FB὎k�*�j6��ҧ	A'�<���sᯏo�Ө�E���_j���(���G0���5����j�i�2���v���gW����B�C�?L�k�<}&�{��JoZ��g�o}ŽƮ��nU(c�� ��g��jv���)?�ï�è��c��Z�u'
����*a��Rz-�i�;|A��.����������w��u�@1��8#������ F��h�w4h�n�3���h?�V���$@ZI�Ƭ���0.q�犣��QY��i,���?��y�+u���L����1[����u���2�ɪ���P�E��������+S^��|=�ƨ��Qi5���V��^$�{���]�<`�V��3�W;�;�n�ww����nT����ޕ�^'֭�җ����������o��T��z(��/�֛�g�_9��r|H�?����Ca�6q�����ON�gߊ�[x�[�8�R{�4v�#~T�����Bk��os�+b1�y6+G�7�s����"�/
�B	�Ƶ�����\�}'𢯦{�V|�[y��c\�m�B�d�.����G�]��5ܚ�R$QŪ��E��I���=����^mLG4��MiQq�4�I~�¬"}m"����F����1�N����$��gIÖ�l9� ��V뜷�$v<
t�g=��<�I��%��}^���+�ץO7��P��p��ib"����P��n1��t�[%��	jS�Ӯu8��i��ˈ�.�F;8P�<�늯���yc�B7�ev����:L���ќ��^��>~�O�Ŧ���^
�r���۝Va�ѡ�s������|#��m!Mf�-�,�R���d���2O�]t���N�K��*�^�:����2����|;ai�^6�br� Z�l<�L�����We�D��b�#wRHl1RI����m���~#���y�mup�|_2��F:�N~F �F+�?gO�z7���Yk��%��u�徙`��;�%�s�#�\`�z�{X%I-L�巪�N7��u��?j��$��ŧ%���
��3�789��>�v
���\gA	yq��.���7�{����Z�������躿��~iQq5���<���s׊g���3xG㮟�M�i:ދ��c�${������?ZӖ��i|��V�S�(�|�m�o���F�e�J�H�ܢ�#�S������et�O@[f��ڶ�$����=^L��rN=�}�g�|Y
���',0c��Tm�L�{~�� ?e�����_-��b9�{�Kɧ�_=�`��R�[}�eUiSr��xͽ��ח�MAd�eRuMY�1X�� <�9��:�2ʹ�k����/�����s��<��;Wq�C�֣��\����dӼj|ɮdS����ُ��`��� ��>(�M�֣*�K�� ��[~i`P��W�����5�(�kT��Eh����]ƪ�7��wb�vm� ������t��.��;�L� پP�]�R��jQ���3�3�OS������5���Z0Ӛ|�t��ڌ�u9� �yz����Y��.Xm$�.�� �����ϕ� g#9=(���G�k���֋���3�>(��n�ȵ�l��U�[��q�'9'�'����w�9��OL���������/�~^\x�@�%�rN����������'8� �?�7�}2_����H�ܶ��:����y���z����#Ω��e[��Sã�����?���o�5"1$h�'V�@�WG�mH��Ά���pc��DE�������_hi߳��/#�{e�O��:���A��p�����p���:����<w�;_��K�?�Zu̍u�=�W�D� �H������gV���c��U[v�yޣ���w�|_��~d�Z��=�	�*3�Ns��h%�_�>h��tj�������/O�+�������|@���bdwr3n�Rq����h���O�������e��l�]1�� v�	=9��J�/C����N��Wř>�T�4���ևmuX��[�>gn�FA��ޱi�ي/5� �?��<A�k���4�5>~�.Iq"�����>,~i�����Q�
%8� V�c��>|C־ x���Kn��>�5ϵ�6���Ѱ�� �G�~�ׇ��;Q��0rT䮙�.��T��[tM�ݹN�'���x��T�Y���ҿB>4~����x���V����lZ�1�ci������O�_������w����~�L���"@6���f3�Wg�SjJ�鬼P�(b��F^?z�֚��h���F��(q������{��Eië%�ÐŻV�����x�YXƲ:J���0Gֱo<i<y@[Vi��	���`���fjz�򁑃�#��b���x�S#2HU���ڪG��d!s�{T� �x��O�uͭ�6V�q�x�;�Dv�&��3������w�62�O�}b� I����,m^DN7�t�V^�2vB�Fk�;��P)����b�Z痶Q�~�/-���5���+���ɢ�D�n�}$�娎��O��c��}��� �>��ƥ/��1�1�ݞOѮ�2@�ϝ ��(r�ܛ�	��k:]���_Ʊ��diziS�㴏��J�c������w���~1���}:�.O�g�\\�� �W�:mׇ|�>�T�:��9��*�e�=�|?}��\�.u-W�-��p�Yn'��I�9�'�t�rT���OS�s,�4o
Z��zM��Η�iQk����%ָ�dw��dV�L�1\���CQ�4������-.�-��4'�q׿Z�`��=5t��!i� f�3M5�*3�!�p3�3Ԛ�������̖�j�����~���NEyќiE���ΫU����S�؏Z�4�ٯ�W��#S�����4�"W		�p#9<{V�Ϗ�@g�-Z�&Eh���m�6R2
�~��2�����?dό��H����Bf]�Yb;��=�ؾ���������؜��C�����N:W�����t�KT�ײ,%,m(Ө�ц�1�W���឵�q�u��\�q���s׊���Դ�O↡&�ዯi�����n�I!A���W�fFE���?tW;O=z���P1�w�F� ��i�#�85��A���T�'���xL�	�u�����-�b|3У���k����.�gg��0Ö��q�?Z��~^"<������/F�S�u$8$n�����?��3��d����W���0��nR1�$w�;���5�Ҳ�Og/�iT�S�'�H�?g� ��|E�+Q��~��+�V�F{�>�+r#,���wJ����g��_[ġb�W�	�`fF �����=6K/�{�����Be�� �q��W˞7�i�^&��-�o�v�Z�D!%�I�_¾��X�%:�����>�jq�5f�<�h�ēHKp�I�i�x��?�Z�m?r�/� ��������Z��ǟ���� ��G]WY�R�na�9�c? ����w�C�ߏ��]�>)�����%�j������BynS���j��|���d,�+�}O�LL�%�$8e�.�W����t�����;� 	����D{��� �ng�k�M�-�.zg����?��[��1�4{�{�>���\�r��6J���~��n���ɿm%����A�#*r~�6�뚪r���ve0�K�]^ə��	�C�.�~2i����ep� ������~�:W�l���⎋}q4Kn��ZB�,jr'2�Y�8�o|
��4� ~�v�xv3�J��B�!!��N���rqU�� �Oky�|W���fa7��m$Y�Q弹1®s�A�Z7ut~�G	��lyW��h~,��v�w��{Tt���]�\�^�S�+�~c�Ǎ ��~�����P񇂴6��c��X�O�ˍ�0ۻ���9�$о
�x�K�\����WZ�ҖK�ʲ\|�4p��"1�'�zׯ��
�� O�^��[\��w�}���\��7�*vn�ֹ)��Nzj�〓�)NZ��~�	����T�,�.�[M2b< @{���u� ���y��!������z���Iؼ��2��<9��5��/�ak�
9t�	���j����ͺB!9��CW���kL���l|!�� d�Pi�����:ŵ���k��]#:�:t$�5s���|�"�
?�'� �����SX���Տ�o�/�*G'W�#�Z��+}���d��F��O�rG��|eD����"�3��z%����8�;���b�����یס��t��P�7Z��:l�+lTl��j.Oz����_s��Y��o�aЌ?�늼�u����6�}>�T�6y���s���K���>K~��P��'�߰�?�N����� r:�<W�?��>�?�����G_G
�޲��*~������
CҖ�"�N|��lkf�^�4U\�5�#�د��������_~اo�{@[��>�ψW�Ϟ��J�۩�P����J�d�����������"iQxV��>(��ֺ���bo��6E�3���݁k�>]2��W:��K
�m< #ix�G�]�|]���qk�����l�2�F7����
5�ٟ��
4eks�c��R�k����I�I+e����x�H��ɜ�c�?͠�x���ñ^����7ʪ�ǒ���Օ���r3�+��)���|�g�;;��&@q��^���Z��<?��k��I��ok{pvƓ�%C�;O�^w$l� R==�+�bf*�$���>��$�����s�g�J��6S��Z�OI
�akcy�ܻ8� .q�X����'�_�3ax#Ǻ6��i�m�D��̠nb��q<���־vk(U�9�'�}����T*3�ۨ�tǥt���=(�R��(Y3�o����;��^��-@�Vp�d�xu37� t��\�K[������h�8�������t?���\Ah&�)��.wg=:~�WG��5�
�S��~0�h�j��� @fM�$�lJ�zW&3��?g	Y�����O�����'M��GT�޵���95��䰖7E1��1A\��<����,|@R�/�����y��_����~�)���|I�;C�3%��WO�@� �n'� �`��x8<�������>�3�e�úQ��Ϟ��)���j^BLV�rdgv>�=j]�Y���#J�����x�� �͒#ν�_��n<J��]��VX��e�'��޹E��|ga���~"xX�D@_I�.:vp}�_Y*�M�I&���Z�h�p����Ce�B[c�����>1i�� ¥�fm�J�l�tHįˁ�=�k�������㦉j͔��>�	��?�o�o�kk��K���Ls�ڄ�dS��?J���rUcS�-t~�. �X��Y��u�e��X��`�V�r�~aS��|A��k[�n�g���+*��lv�k�?����� ����W_���SE�����'`�7aA�;{�����|I���KRq�md� zW�⩺����?5�ƥHK�]R|,��iq�Mh:}���//�иyTas�|���=MyůXk_��.��I[�"���,r1�1ڼ���������h�_e63	b|�=s�Wa�����PTE��s� ׬�JqP��<�ك�AA[C���|7i�Ŧx��᭭^I���RX��Qd|����V<)�g�ڭ�K�S���D����QG�E9�������C����Ku-����B��9݌rx=�W[࿃�$�ׯn|/�ìil�^�Y�q�'��q�[76��� �˕'��c�?�-?��g�uK!2F׆G�#��sQi�^��D�|y���;��#�i.mI���ԃׯ�+�Ծ	|X��8�-&���1ƾ\6��2H���s��Y������~"|@�4KwU*֗-%�����+�����N5$ߴ}�k�ZC�kZ����ܚ�*:��A$t����8�m��th|�O[E�������O[�0'[iC �G�y������z����n|y!��B���Xq\q哺f����W7�o��[�u�-��׎G��Q�ϋǄt��DռO�]?�&���0!�1��<{��O���\��ǎ���`��ߪ2xU��i�tW=�� �u�9(���eV���u��>#�u���C�4M?C�Ok�i�R-�0�K�bI `���=���M#x���x���&��� HM֋���A��=1޼W�wx���;F� ��k�X�n<t2*�� �֪�֊GD1��n�Gs�o�0�n���o	/|��D�� ($� ��M���O�#����B�+�D�6s�˷�g�+�>Xe]��<B6�eP{95�tK���~��?���e	u丒5�Aq��=�7'�"5��-��K)��L:�ԨZSx>5pA �;G>������*�_�6X+�>���}�ֱ����h���R���_�r�PI�� Y�db��@{���wħ\�#첹�ԗ�ׯz|��ΩKȿoyEu;��p҇[V�]�X/��zVL:���;F|N	%�� e[����g��/0�95��q�A�*��<������MtRK�F�H�1���+�0������F������$������ �MC6����� 	39ݥ����� �pB�<t;���� ~�� ���D�����[}�'��6����)ml���j�m��S��;kl��.N����ַV�m=�/�VO���6M���i���=kF
C�m����kȑ$�C�2T����N�{���0����i:.����M(�{է���l�5������f��Iu,t�<�2��8���:U�K�#�c�:��x�P�#�Q��p8&�/����B�e�Gη��VK�{�{c�G��5&H�t���w��t�c�ϔv?Qڦ���^���\��W�Q��0c� �{H��%1�����7�v��~����iV�� X�_m��D;�$��?fO�z���}�Q֯E�m�wId�mQ�q�`��U����<��j�E�t��5).����V̲8� �{���F��>����S���o~֚M���|2ӵ���Q�,�tl���� �����/[��
�c��v��f[���g����=+Ϳj�,�-'�-��]y&���c�(�w�\`~u��d�`����_M�n�4����5�ĐG$1"�˶�>��u�����RnT�Ij�T�=�/�
_�����k)�̳I*n��8��?���\������4-";�{+=Z4��&4B���Nx�����ȟ|E�3�Z����I|G6�_����'� udQ��j� ]%��_�*�w75x��̄,_�<&Fc��Q
��SEBP��/���Yi�k3��9����@m�i	�_q|Iy�����մ�.f���$��w�7�B`0�'�@j����Q/���RF��y�ت��'�$}A����j��6����j���/�?�J�t��A!�A��ް� ��-�*1���۟5�_�s�w��/ci�=2�j�ZD��Lq���i�9۞��1���xW�τu�7Ɨ�:��:��_��PN��UY~�:�d��>=x����1����
��76*Ybh�(�������ړ���/B��5�!������ R�fr2\�N09�l����G�,US�6�~�m�]x{����l�RG������l��+�I��72�Ğ�K����|w�{��׊tR����$D��.<��ڸ*
��q��Q��?/>8~���-�]%φ�ɸ��4��nn}F1���?�'|����'�Y����jB�'�h@ �A�'��]�t8*T�]JS��B��`���%xF��w�ZO�}v�k8�,�6�+�c�-���5�W��X|c��%�6��� f�v�2�� ��ٙ��u�s�G��n�$�6���h�_➝��m97P,+q���1���t�E�O�?�K��mi�G����jL�4:U�t�2Ȅ� �nNO�^��U�Ź�\y$�m���|s�KǨ�Ɨ�`��E���j��ʎ�=}Mc����/���z�����+�^���X����]���rA#rEz�_��uO�zoÓ*y��V$x����C���Z���|7��ko�#�.�>k9#��TJ�r��`�Τ ���qb!Jt$�9/&|��7��}Z�-Z�V��Y�nZœ�frf�WG��/���]-<�]ϯ���lnux�XV�m�q��;�[��:m�����}&�
�qr���7gi#��#�+g��-Ѭu����G�y��-��<�ԹS�ߟZ�RW�X�~���{��W�R�>8�3�]7MMJ��+��A�T�Q���22�3ֽǺ��'�� �,У�ӵK+��ҢH�{ɲ$x�7c=�Z����X���x��1��hZ��%�-d�h�P�)��$�sޱ�W5׌�i�	i^�jsx^>�T�-�xmR�ď$g�Z�z��W&�7>�V6�)�վ6�w�__��l��|?���f���m�1�*�һ�c��S�߶���J�;𾝭hwHL��ǆ�q$��#8\�Z�� i�k�?�kۻ,��L���țmv�k�dc�OR+�.��ʛP�iN��d#���fbx�(0aְ�^�j;;���fX�uڌ���^2��?g���|�5�}�߹T�Nx9^�ꤎ>��� � �O�U�����4@�	�sc'���&�u˭.�wQ�O�]&��O��N^�i��?�mi>%����3�3���J�Z�c�H�\q�����]4�R�H�(�4��uG'������%�}�WS� g�'���s�'� ��]Z�P���[\�FVW�t��܃���8����E|koYj�k׺�M<���B��W�� �s֥���>/�� �-��r�o���kP�*W���[}f���tmw�M���Ɵg��~���KX�0}��T�A����q�+M&�����"�^.f�0�
I�5����#]�:?�~"����4�Z�$�H.7|�p�ݐyn��׶>���s��N�g{��n��<�߆��[��T�1�=2���5�E,����q����O�'¾�W�Ð\x�� Hp��ق�l��Z6FY�*1��~]���ǟgMP�
�sCC�Ӊ���gȐ���
z�m拨iWPj�G��f]�2���$a��'��+��)���Vе%c�������ɹ��:���Ó�pF2C
�狕M��e^����q�#o�:��_��<-�4�z���E�y �T�f�qۚ�o�\�3^���@8�q�+�񆡣�g�E�6m`FXk�\�~� ]����� g�վ�ˡk�Hm��r�Q������\���nM�3��o�����'�t	�eI�1��g�rW��9#�W�B58ṓJ�������tfT �:W]o��V�K{Ge$�Ȣ�W���]�wNث��4����w��.����t�>̝���8��֦)�^ǟ*j���z� ���� �jQ3B9XȤg�7ϯL��'�� �ÿ>��wP��+˻_0�a�6���:�MC������3�Z����kG�o� 1�{6�d`��z��QO���xQ��m4���MѺv��O����Q��m��˱�N�JSI���C�d|>�����[�cq�0v� �^O9�J���������zQi�n-�7,�de�$v`׽��_~���҈ۂ� ���h$���ϡ�1�����.��.4(.��l&�	�\eB�� t��|׍K$����ԥ�ќf��V���7���~�k��K����}}ydI4��r�3]t�P?�1���C9R��<m���5��� ���o�*�E�~�%��H��0��Jқ���?��# 0pN�l�#�+*�_^n�߼�;0��jt�Y+$P��~2X|`��|E�i&�ʹrS�ǝ�4js�C�|��{����c��i3��p�����$8=Gc�⾮�k����]i��M�u#}��*H�pY=���-���|Dt�紸�{�ay��+1;���+�T�a�-TO�̳:�o+˚���>�#����^+�\:�k�%��ؒ�A�Fl��h������ן]�W�]��o�x�V�vZ�Xi��8�%o�H� ?�x��>"|f�~#G��M�i�N�� X@����}b�HВ��Ā����Ou�Q��X�4�CU�揨I����Tq�l��A0�\zWdq$ށ����K��>9|i��G�?�s�M׌w�[���IHV9�݋��|��e��ŴK��'wI�B�1'����_>%��3RMVm�K�>f���v�� ��쿲�i~$�k��:�v����U�RX�P����iԌ�4��1��!W'��������� ������Mo̗O���_3Ȏ �$�nlRA�����_��ퟦ|V���=4�됝�ֈ�y�ڊcf8`�<�U�`?��Ig��3�J%�[� ޏ���89��Z����-�>+�|A-��@.[ɶ�v'"Gd~X���5�>x��\��*ӲkOT|�῎PxK���ݽ�����\}�`��m��m#s����?4�?Ǿ�Y���z-���z�wE�}̬�O�T���a��'�O���|_����p=�Ѽ�~����S��;ьd���@�����⇃�T��l�5�`�˫=̑�!�80^F:QEIK��#�ޤ��s������������u�=A���nՄ/|2��c�5�_<)��w�
w�}��R^�wIH$c'֭��G��݆�� ����ؖv1B���.������+���'x[�_�S�V~;�%�����_�c$�����o�94�9��j�$����ߴ
������6k�y��b��k�^���]N�[�}�;�e#pr��f�3�߇t+� ��3�����&�,�L	)Rr�FXu�xt��O�P���k{��?(��e����#�k���ܣm�1�q��C�"�W����J_G��!'�@��=�i� |K'�.-|7v�.��%�͍�d�F����Ǯ1�2kx��}�����,����[#�}���� �-��e�Y�����Y�%v���<1�⇻���C��7:��v�Pc�X�+v ������Ȼx�G�X�w���u1�4�)wnK�J�˵x��X'f��<J�Q���V���b�G:N�I�_�ҨG�;V������|��忠��M�cJ;������*	0I� ����J�;�|����~C���_�+����-���S��O�uQV{M�*u4����_�k��)G�,{C��>/���S��W�_�fW�E��t���d�͈қ>g?� t^����~���AE�U�э�6�N�};V���n���GoaY[wK���c+���*E��aq߁L.D�t�4�� Y���0�2��-51����e��pi����2��ȿ9��P6��zT�;w&��W`�G�pہ��}�K<�hU۴���� �_ʳ��+��}֡��HL:ִ,.�]�� g��+dn���U_�Im��m����9�<u��HX�ƺrI��*�й�J��~ƿ>�g� 4A�������c���q���g�eyU|57ky�:C�xh%��e��p����g�ڸ�o���t�];\k�Z��h`�A�Jwb��� �9�[V��Ԁ�0/�A��|�~��)������^���	���s�Y�}�~,���:Ӵ��I��&���ҫ<�} ��ٮ���^��Ai�]_366��W�~���� ����J���*9�c��/
�����o���S[:�֒|����g�'ǞXK4�j��Y~�z���঍K���*�L�u�� ���L��~X��n'= ���+Z|�o��Z�U�sErZf'X�Ҵ���bQ�v1��鿉}�}����.>�y��O�C�qR/ů�����	�����~��>x����7d���z�4� ��ᔒ��O��~_��������g�`b�}�N���.�G�_}����I���P�:���|D�/�C��d���I#q.��׷n��z՜6>"խ-�ʂ��H�Vb�(|� �i����8��r:�ʽ�(��J3�ڊW�j%x�8O
��M���yjڍ��gK[��݌f��z}��/�}w[2��D�Z4H��s\�%��@��ֺ/�������� g��zv���6��y�B�~_B}k�%QYnx��ڧ������W�f�4~� c�����1�F1�4����5��՘#Ɇ��O-̙ �8���g��kV�Ek�p�"���0� I!Wh$��>��ǧ�|�`��%�t6ŋ��=Y�8���"��-�=�U�[���!��ż�$��mBeV��_d��< @#,pz���Z_\Ay��'�w6r���{�?�@�x�/��0�b�x��N׷��d���bZy;<��O�big��Kq}&�5��ykˑ;$�Þ������G\e(.Yu:ٴ�M~V�}����[����6�����X�8λ(�������Օѷ�L׵u�B�욃�%a�*��}ֳ�7�3!�ư�N��UqU-�HGE+�r����*�?Ո�F�/����r�������w�k���^ ������?���К�<w��,��3������8����T.H>�X���W���#-rR돡�ym�C�jQD���+�a�^��b��Ҹ�X�#��H�?�Ub�ˬ��������(|+��-.�Ӽv�&I�ZH�8�wd
~��6�(]jw7�/���/��0�h֮T�����?�>��ň��x�R���5��bGG9ǧ�9�G�7Æ��$���m|�����rMO�|d�eq����<J��5��e����JJS����ڐ�]?]��O�?�PT��q�U8t�]�d��6:��쟯=k.?�_��-�x�ܻ6�ڸ�ޛ��T-|[��w��ȋ�� �P�}�O_j��}�.�����gjrL�_j��� ���mU�p_�<g�u�\���������2x��U� �&�Drm_�Ѡ)Ԙ���KD�%���D�^��CxU��_8��I��� aݛ�o
i��5MZK�u<���y��99�u�@x��$�Y�8� ����o�BK�c����yr4�z�D����8��;S�uqy%���R��ߡj7~���4��/�̼�$��P��,Gb01�5͍�7�$Wq�x�P̚���G��랈ݱ�]��u�mR��]|Gԣ�5V��l$tc�9���[O��D�-�/�?�bm[^RD�����YrH���YI�do��η��ƛ���S�h�]x)��׎Y�Y�t=Ձ�v� ��~�?�U��i,�Ֆ�� �=t���Ā2��ھSկ�~��j�Z�ک����#<� d���W]2��P��+��){��A].�9!O?_ʺ�b'MY�sN*�e�=����A��M���������oD��Ԓ�y�֪��-�a�?Z������R�"�4ɴO�h�|����J���F�s�y}�����2�u+��x�o>l�� X�ʧ��s�y猼A���y��,�"Ֆx�_�� U�O֭T�Y�Q���Zq�3�����ֿ��ǒ��Z�h�@ֿ�P��J�S���j�<�r�~����/�<A2��٤���E��\g ���� ���5�����v���Eo$�2Z��T)����שI��-�i�&���3���Ƽyq4�B+c�9>k��ƥ9���L�`ZW]c�Y�!�#�~_�ڑ�0xȍ���b8��c����7���g����ݏ���=~�H��O��gE�S�e��?-��."�=]=I|)�99�����_�cy�ᎁ�+�,$��)�����F�6�A���5�
>"�|(���x�����r~�/"�*�����:o؟�}�e�ɩH�����?٪K�|3
��jY?��� ����F}��e�iƣ��>q���Kj� �,��9Ѣ��7zU�pX�{���K.A.A� �q�?���k��H�$�,��!#v���d�}3ZS�ʟ��*�W�����YAYM�<�'��
�n�W��߹��� ֊+T�;#ù�&�:��y����\�ۢN�G��9����6v�
�C�W�r_?h�c�F�4p�uo]8{�!�ۖ+"I�U����}9g�%�1�T�4�Cd�#7�+�� ���G�>���v^���+�I��M9����=o��b�(SVg��d��<eI-;���ڷ>������i�95t�[ ���z�_5k5��K&�����G�c�,n	H���j�N쁓�#'ڷ4��7��>(��lw�W�!<9[��d
!1�YN\s�W7Źdic_�u`�yk%�]y |��@O5�N�ih�>Z�6�hZ����|F�4���7���q���fva�s��	t�އ{~|9g��E���=�D�ؐ6���ڹ���4�'O�7�$�w�K���� ���|B��%�!��%��څ�D:`PK�W$n+���f�<;�TZ�܆��k��}"�-/�,jQ�R�B�v�!��A�8�R����o�͠�q&��ݬ�.a{�Ky�:��8��ω?,o4�<-�K��湚��u��;�b9#>���8G�*]I�+�R�����jP�lޮ%J�,z�-���\Z�wڝ��͢�]�nF*�6���x�Y��p�����|l�ߴ%���P@.Nhk�#o����i�z�/�Aַ���Ԡ� ��g���)���3@��t�Y�Ы3�_r�8��]4�5�x��'')�_�����kM�{�#�M[i<�p��� ������j��J��|+ag��[/���oD8Q�\7����pay$힟�H!_/n�o�]I�s�x�S�{�>4��c����f���%�;�}˴�C�>��^�&���kW��sj7V����/!q$��Yp�[� g���e�v����H!�1߷�*9���es���7��K�Ѽ3}w����������B�}0z�R;]/�� �Iy���wMa�Y6��� )Qo(9�8�� ��8�|��2 ����*��	2���@o����5c���sO���i2�KtI|C�F�����f���#<7͵�&�����J�u%]i�_�O.=B<ǵ�G�	�~`��>�������oŎ�jv�� ���60!���F��d`xc]'�4u�:��dR&-.���[�7s��2��s�~����R�.V��R�h{Zl�X���b���n�[W𮨅E����I�T����j��oU�_�Z0/���?����.�nnV���]�sl�����Lcy����Vy��5[KҬ�R��>jW)�"Az�A�C���Toˡ�Zlׇ�z�ڔj�
��Q�߲���؎6��ڬ��#P�5�]W���ep����z��i�Q�V;h��SSk�\{E��_=T��x>�gڭ���[ƛ]����ФSI��d�m�NǊ�v�sx�I]�z��/�:�o�_x��<^�th����4�]�ȣB�s떫�;���E��i��&���i,�P/�b͂6���׌w�o�^)���O�>7�F���I�K�ῃO�P,n�&;�7m�J�	�5�p~�� �.5=F���
Ej�R�ko-���9�@G-�8�"��4��n�SN�T�=�	�w�<k�h^�=�x�H�-��]�Rs(gl7�ۜ��ߎ��F��oW�.�l�-ݹ�]?S�RCH��|���N}�5o|E��>+G��#Y�u����W��Og��\��0q�]����j|=���>���o�Ʊc���Iמ2@qӵ*��/6g���J\�4pZ��jZ�xg� E��vEspB,�빎G�y�2wum&�OU�t���}�⸭7R����[��]zSN�d�6 �2��t>�v�x7S��o���ǉ�k+6��i.C��8`I9S�8��)S�VL��!Q{Du2[��YM�GQ�+n?
�&��f�O�ُ
�Q��ARA�S���E-�8$�ỂpEy����W��m"�2[��B�(��r��\�����#	�Uj*}^�����jJ#�մ�z�k�����|;�5�>=>�M�1�WP�`��[�1^�s� ��
�i��� `NJW���D߰'�d�b:�Ȓ_�F
����"���l$��ջ�C��+hyΟ�[ԣ�k9�����_�+t#�.)5O��%�l���1E�=Rܹ���Oz�Y?��_y��ZF�@��?��[�	��(�,�"�� ����V����:�I������yF���5��կ,�v�����nq��<(ۃ����H�s_D����j��5FS�jf�5_�����[ĺ��p��~Tka���t.�[\�O3�W��$����2v�� �Dޘ9ǵD�	|"�� #
�������F��X�Wmjz����.��m��O��~jB�ۺ����<������{���f�uR��O0��i*�	�.��<I���N��|$��bK�0ܱ�F�L�ξ���
�"B�=_R�l[�H�=�_)� �����m��U�	�Qqu#8�2Et�*X۪Rw]�4˱ydT�KCm��я�^6�nL�	U�ܣr玼q�Q/��[�� �Ig����}��ַlu-�� d$�ֵ��R��i�]Mc�yr���s�1�מ��|F֮���9���$Z=�P��1f*['�A�O񯠡�6���S�sͶ��m�� N���.�,142\8i>��6��9�pŦ��ڥ�����]��+7�<,ω n<���?�v����8A\�w�nh�&m��_��
-rO�	��U��v��I�` �G�VlTI��wm͸��S�қ��X��uuu�K�F�d$|�����Ҋq��.cɭ�{���c�Jҵem�� ,[����XPB�f;T �x�j�C�5��ϒ�iRj�p��;3���g���� _�� ��ѩ�W�_��?�M�A��� �_F�}~~����EU�SZ�HzPd��ȯ�� lӻ�=�8Ɵ�����n����߶r���dz�O�� FIXb?�ϗ�l"�G�j�oN3��+$L>�@�B_*�2��W��VF�n��&�n+s�*�ԛv�����-08��"ɺ���ϥE!�0�I�ǜt�8�D��&x4��e�q�R��̧�]B�č0�8'�Jp���T1�?�/�ZE��g$���G�#��L�&?���K2����.�S%���+�O�;�m�������1�Ӭp�O��c��^qnjk�����z2+L��r������d�ܩ��sS7�6|�w�,ɝ��C���x^�MX�m�sI������5���d�N�>�f��Gpэ˷�H�W�č/�G��׵I�1����/s6>TQߜV£��Ov�:��� i/��|!��tݗ-������}8�zc������5	>#���t�����u6F��G(:.z�5�|4��L|\��� M3XY�s��%���˳��1���_s�إ��ii���5����  �`c�sֽ�EXe�����f4ҩ.il\�e���g3X�l�Hd? \�y���lc�����?�\�����(�R�\)I�D�@o�~�z��i�֮O�v��{`+���M+?��ݏ��zE_j�@̿�2��q� -z�?���5������=׊�+�]�� ��ßi�z� �`���Χ�X9� �/�����؛�z��� �9�6��*T��aj�H�(T$�E
�ݤy�Ve�PY� ^���b�t�'ঊ<E�!� �f�v����G��K��׷PGl׫Z�&�s���Yb'w�L�w��-�y���oc��,w�5�^�xQY�>��j|i�0׷WO��i��ԟ�q�z~UCТX�>"x�U�9�����ݷ`���:�+���u�_��m��pv�Q�Em�H_R�u�!��nO��W�6�� �H�l����,����T���]Hv�i��0;T�-�b�K������%e]�]�B�����I�A��k��˥��K7Cx�����F=+{þ��ziHȚ�Tu�u$�}1M�/y�V��ū��~����J�wgo�j��iw>��*�ؼ:��,8�&�O�EGsx<�)c��ڪ�4�B��1\�r|�Mz����x��h؍��Ϻ��*8��<�?�:ylc�*��_/��B�J�@�L�ry����Ѩ��e����s��
i#�������+u�P�(b8by��8e�.���� �_[��L����������ź��T0���.][B����>ι���UhٖF�V/�-<+b���Y� ��P�ÜQҧ��Dʧ��U�[���l����VEO���w��</��ڼ��~_������v����n!Q3���Ǟ��Z^����W:�����VK�\ݻ���i'������:�ãxr9,�+���et�$��,�߰<�����j6L��JR�Ӻ����!�D��8�M5��3�L�U/�L|�� �� �e/?L�Z�O������� ��x~�-�b[� �r;U�>1x��Z���m2�v	oaob����#$��Y^��6�J����9�|�Ԏ��r�[��=���Oi�Ei��'���rH���^@�.F�N:�I�o!���##��t\�y�Si�9������G�=�m��لȧ�YGF�u��Æ�O͉��ȳ��ح��im�<���>%��K˕'tH.	$Չ
˚�zW�/N����:J�-�9���v�+�NHr:c9��Ҥ���5{��=b��w��R��`�'v�x'�O5���6�aԾ �p}��Kf+m�C����6�H�'9=i��W7Q�2��-�J/�o|q��\�A�ۑ��ʇ����t���/��9��o}R�+�`��ڪx���G��7w�� N����5�~L��2)?*�=��W)�eo�?k � ?u�*��ғ0�+I�t��W���#ɋ-"� #�b;x�����k���֚�˽2�?"�9#�� 0��<�Yڡ�Fln;���fx��O�o|�K���s��U(�c��߼JG�?����Y��u)�y�>k�D��'����� �y���U�jL��{�|a_����;~5��ah��s�g)I`(۪��
�w���9�h�U�z�zq�l|�*rvH��x8ە����<��=mEm�o���Gj��5+]4�eb���s^���Ձ�d���*�w����]OQ�[KG2?�=p�;����i�D�i���*�-x��-},ҫyV�3�#����Ol{����3�{���"�����}byɼ	��� �{�qڲ|u�C�?�Yc�C+�ټ��a#|�����'$/��}w��hпg[h/��^#��ڑs{�4V[��9��Ǔ���ʎ[j�sv<�ԕi�;��O]|<������c	yl63��_���|��~ڋx6>X5���	�ßξ��u�U$�Fe�9� _"~ޒ)�ׂ��b����?��^N[8�Ʃ�x<H��]U���E���'U��屁S����W8�
�VlW�ڤq� ��9�+�)�u��Wr���z+j6�<#�G��#x�Y��}"����s��j��Qo�ZF���#1v䟑�S�EU���LA?�(���v��'�w���q�6�j�ZNI��'6����� N��F|�	#���n��Y�߄�����l}� �\���x1ϛ'��t�)� �T;r��ޕu����1>$���0���U �$�;�z�qc�sK��u�N�]�%4�@�#�"s������'��,/ kk�v�$M�O���j�T��g:�����K�3֤��F����UN+�ɟ9)(y�S���R�zf��6�.g�@!=�DS�<�*Ì�[h��-�!�!�q�>�#��ץ|=��jP���x-n���#Z`��c�)��#p9��ǜ�d�N;b�\Dh ��9SU��=\.*TZ]j�!�և�N5����Z�<�t��Kyf'�x�� #��X���kI<?�e��<�E�&9��9NqU<+�;�Z]��|[��|�/VU[v鱏u9����_��l�Y�����G�8�wԀ+��]=Ϧ��P��`�;��� <��<s�]����k�����p��9�}�*��~+],�v~4�����3q���4�٣c��=���.n���V�F���b�Q�ʐ2��A�ҸU`�6����y�s�ְW���u���E�:��w?<Qe�j�X�Ss�j�2�rm�����s�ns]F����~0���ĺ��!Ѯȴ���Uc�2ܖ[���x��4� & {�x�E���Z����9Qנ�&�*�A�κ��O�? 5ׇ�j6�]��[�	a'���
��0 c�N��^��ޣ��O�_N�4�3��$;�,OZ��� �Y���ܿ���|�3���ƝI7F-�,MZ��NR��f�tLG������|T����·W<�/��69�>�Z�$�a*G~��pz���W� �/��t����K'u9h]����vǓi���k��8�CÒ�h�K�l�̵�.� "�����r+� h}��?�������[��ezci�������O��Z�j��o�q�5f�GC0�$��S����)����+�����n:�I9l�m�x�j����$o���GJeΤ�B����wt5�x�Ƒ[ö2�_���+5=�
Wz����c��$ �lc޼�R֮|Ap3�/�6z���p�Fl�
���M3��MC^e�����W?(:�]�0��OsYT�8��z����KK�DI=����1�����OS^�Z������|7���,������)m�`�e���� �l|=�g���G\���y�+�Q�#�$��V��t=�5�G��/��5�@𶞺v�
�y�c���� 5�U���աg3�s�-�'b�4����Z~�����Ad"��)�3�b3���o�u� ��V9���_��l�J�%�cdm�q��/��� 	���H��>��j\Ҫ��r�sN��%��t�.Ӹ����*b�0�p3��s۾k�ev��]ǟθo�
�����������a�6��������3�r����S�;ķJ��'�w�3:���
Tϟ��O�$g�zO��'�UG���'ckKr<��`� ~����j��:S�������NM�B�j��)]t���|�H%��m��{&�=ML��pw�ֱ�"�����z^�Yr|� �q��K�i���}���߃g���O���r����G��z��?�����
?tʿ�����*�X)�-#t�79�Wğ�z�������?��_m�O�&�)����\;������Ez���-�6��o�<cXU�I���*�Q�$�z�Օ��*�3���?Z���;T����Kp�6�3O#��}rz��FM�#�R��Y�I����1�U�~m߅u���D�+a�ir�d�{`z��8������2/9�[aϝ !3�'��Wi��*Xg{o�#���H��[c�`� Z��>l�}�{����i!$�~@�RGnwc�åG$���@���6�}��H���a�	s;0P���U���!k8��HQCG ,F	'�ӧz�b���վˣ�|7���X�E�mF�9]�OO�X`��Ҿ �������X�����\F5	,�,��; ���E�At]:�x|)�k��Bo�|uc��W~',���\���|3��Q�d~�\|l�M�����!���	Ķ@P�� q�sָC���t�%C�˯7#�h����q������GĚ�յ�Eӫ���"�	�t��x��O�MZ�����C��J7g��1�\��hGd}uOim*�f� �w[�B�i���Wᙵ��(X�+�;��_��_○����,-vm�m]�E�;�~�c�c�>;�C4^Ҽ�-��j� �(�X/��S�Q���φ�Z=�>�u�mf�����\���K B�$|�dt��r�Ys�VqB�Y{�g��~ɾ:?�uMj��-b+�%t��x�\��>t��C��A``s��!kiuh#�����1`�X�� s� ,� �kġ�ˠh�SǨxR��a�m`� ����$V���C�J;8�.|�+l�Hl"�������e�q5�S���a���X�f{���[�kK��W�����A-��^+��#�#?�&��X?�o��S�U��R�ycv�v��2���z^ߴO�.�R��<�v즎N�{��_���egmr�]���Q^�F,d�g�_�x~^UN�ڮԋ�1
��I�x�R��I#���Y�I���$C�{/ĜE����q��%y�ğ�'�:�����@�Z|��F֯n���
U�H#����>(�� �w>N�G[��~ux�S�$<�X_�ׯ
��S��G�[xKKּf�tz���PYA1�F<199���\g��A}�Z� Y�.E���4�:p��B��POJ����� ����y�[�XE-̱#�uC�q��z⴯��
�VU�w���PI�޺��Τe��MI^�5:O���}��󄊺T�'����U����"�#���0ܣ��O_J�����E]WO�h��v�9U��<pFO�T>��Ð�]���m�c�Nra����:���#)a얦u'n�$'�H�ok~X%���oBd>�O�]t��B�L����g���?�/,e��L�������ޅ�y�q�W�����t�.�s�oo��Z��e]*��ɖ�m�8�H��\�c��b�A�)�:�*94	�w�r;�y|���~R�d?�L�!���|���� v���7(皸�X�N�጖<�=�0V���K��+�Օ�wd�sH�Xط���q$��]�(���9 �z��z�^�㧌�ѩ]Zxw��ta�a+���8﹎~��t�<���%�Ke���O�<̹�S����+������H��SN.<G�|yڨtO99���]xx�S涧���)E6����
�Z���ǅ�N����#۶K�^�I�=���#n��?�)a� 	w�nO��#���q�U3�xy�D���⁠y��0��Q�����G^p=k��\:o��"��u���9��0�q�`�$��{�EiKH�S�RR����5O�*�-��49�,4��Ձs��b'���{��#iZ5��x��?�/�*�X�3�pNX���+��w���!�i*H�`��I۞�5G�:,z^�/!:�R-t����+��f�ӕ-R���e��ox�/�5�gg�u&��͋��'�z��-ż3�O�H<u���D߿��	�g�L�|�����z����&�>����S �H�$� �9#��k�ծ�O�_'�ʥ��� �$M��c� 7��mT��X�T�z��g�/�4���}Vc��C���Y(?g��a�9�r�I\pN�\_��f־+Y�]��\\	�I$o����z�{S���M�4t�t��iQ�g"Iʺ�v�$��#���͞�	�m��)�f��5�Y�2�p@_n(w�&��n��Wc��|��R6�v��
����6�*�p9���+��,z��ZLf��|�vs��9 ���B+���60�FO5�����>O;����Nj�_�[�焒�9�����I�Լ��}�&�m3L~�<nQp� � ����)���!��X�w]�*��PI!O'��qV~��[�+���%�B~�m/�s݉}����9�G����3j:�:@��D��bDV������=k
4�^jh҆�8�F͟Y���:��~�iV���#k��Y��-�2�,�=P�K���r�wR�^x:&#�>"��z�*���<E�G��L�|Nu��;���x��������ſ
�����'�q���}���Z�&9T�O�\._W��8�Zwj� ���g�� �@��r"֡m����\�������:y��-R&)�~Q�|��κ�~q�K(��B]a$c샟�5�����ۮ-�&n]���V �=�9�<?�n܁UV����������?��=X$ڈ}����k��!|C�_�mr��O�7��ݪ6#���m�w@1�^%���X⻾�Á�#�o�u��`���{�9,0_��دY�E����z;�Z����ܮnS�����8��N��a�Q�p�J�5+����,���u�4� يO_���x�_���g������f� �5r�p�{׭�������R���f�?{��^kg�_�0�Q��
1���_��'?�[_�_�e�S����� �6^�rG������^f+.����Ջ=x�2������I����F�Y��D0�$��O�G�W�~�?�o�ڧ���3S�&���f�R��pT����=F�/��0F�h��l�O�$ӥ]��/���3ľ�e�|ie�i-4�{��f[�q�
:�c�F,�B��ٟ3ęn&8
��x�:b �<���3��7e'�#�=Ag�=�GG��_�-4�b�f;�@,F��3��Ҿ�_���OZ�O]M�d-���GͣG�9���Q�ğ��(29$���<q��k���N�x·n��%�H�3�u�'�d|3[]"�x���ae:�n�!"W �'��y�������[�P�C��x����ϓ9�����_X9��� z��V�4�t}Qn-�i�U��$�9�9��]Ο�ؿ�� �t�ź�1��O��e۔P��9���f��z����6%~�j��:̙�{�a�`g�6�$4c����\���h����$��ن��-��;�]7�;X5+�<Ai1�.�JX���� q��𫩭e>�����s��}*A�O��c��z���50 /�]os�d��Δ#ބ��n�����+�
탌T1C-�]�M4��,c&��19p�Ck���K��|8���3ιu�D���@�q�;����=����I<޷���m�ږ��h��Y�l��H�/�U�����*��c��������6��6�uz�U�!�bA�j���d:����t�U���A�#(a�����ZR��h{|A�3�yR�2ctd� ���r>�pó��+g���ׂ�����:�qU|�Yꚼ�z��[�����E�c�a������KO���?Y]���I��8�N�q�mܩ�T�R�y�僔z�|7e:?�W8s�6�C�~���
�.:�<Wy�ht�'D�u���5�*�mL�� ���ErW���t_<<�z�������8�Z�Ҥ�Z)ѥc���D���p�٦���Y*�8��$d�F��<V牭��K�q�W}���DRH� +�|8�����|^ͬ]ܼZKy�.Ii7|�ېFJ�'RLs�u��B���p��:��d�z��?�mx.8ǀ|m�7yP�F5���8�� ��&i-uFi�o��Շ��ֶ|5����tk��#��HW��1��;��U(�P��6�&S{3���z]Őp����z�ߵm�E�?�i{���1������� �Z�F�!�@p �3�ďz�"i�WZ�خ�Uѣ���$��rs߂+j�����o��e���G�C��r���xX]_|w�_N��[�+�g[M?<��fؤ�H �5׌�|C����t���v�#4cU8�7�@dg��\Em��{}~�HA���%\�t���q���8ui�u>�%�����i[]O�/nO�����sc�v�(���$�H�w���?n�M�F��"�b��o�e|c��}Y�m5'ԥ���d��:f����2It���%K^�!�c�gڼ�
:�(���Ek_����TFt-aQ�4@�U�o�Vxb�h�������p��4���¼�-	�r�W7�����I�]�1Z�隵���?h3E�MBE�8#��A�q��`�k���c4p�������l�G�S�I�����\h��
��K���*��}��^�K�[^��)-/m���d�h@��q���1�N:V�ï�4Z���9���]}�T���d#sr@���>�B�+�3h�N�NT�'���m,%]:q����<=\4�$��Lпk��z��a�� �{KX��Ν)���A.$�O��
���Rn;[q`�Z�?�Z�7�4�J� �P���[�Ҽ��)��_;[$�ԛ����J�]��IV��=C��7��I�7J�׋�g�9�m�,Ҁ�d,޼��Ş �^�ǚ�Q�%o8�re]�l�a;N{��>��*^x?�:}��o�m��� �Xu
��zW��� RM�Z^��,��ҳ\�O��I.�,��,�	$�G,�a�r�)�6~yƘ_���4����5��p�K#6c�S���J��,�X�����u	�(VAh��>�����һO|d����/e���C%�d���`� �;��υ
m�[y5�_���4���>#�8 ���S���G���۽>��a��9�(��/
�7c��֫|l��� s�����T� ��<q�'H����yp�.�&����ٽ=1V~7Z��N�0���P���� ���[�T�ov��r�t������sRG�G�kh:�x/D����6���`c'�kKG�y�k��.�j��y�y�أ�?5b��%c��IŤr��95�cn��wù����4{�x|�)���{��-6�twe�,J��:��Ѥ�1q�j$]uX��מ����t�(�S�.��]������t�t��nD�;F�F6�w����k�����Ϲ?���Č?�}����u��I<�8�E�ɏ*��dFms�y�Z����.�A�%��{"jf	A:Ť*��a$���:𴌈KھP�������`�im߂3��؁���V���6 �eQ�n���C$y�DGvk��Q����WM�\��w8,@*��~�YD.( �m ������}Zzw��k�z\����)bph>�*�kC��G�BǗ�(m��������xE�uN�C�U�j�ysS�C���V��W)��TaÂ�.����R�b��&�)�	�I��V���R-B
���W�ǜ\����T�� �h���p�6�Ǎ��{�~0_�k��T�[B/^��\Q␲YC�ܚ5P���ͣ3�^�F���V�ZD�Aj�(?�kn����ƹ���T�O�N��s���'n%��[&��ͅ��rѮpt� %4�i�seރ`KB�^S�������)Z�JID�֚J���`Y�	�O�A�=��a��.��i���p��/jq+FbP���.��2�>�fʝ�D|���C��%�-��?%׿�'��n��PMIkd1��˒�h�'��-:){�&�sس���{~@+U5L��p}��∦������Rx�`�� �l���<�h��<��!�u�&��U�z�KxD�.���h-a6�6�`��_�
i;@g�����'�TXh��$y�l;p-��G0Gy�D��8�n4�`�A��V�(���a����L�Cs'��X�D��$C��L8�X	L����Y3VV&`��e�8�Tu�h��<4��P�@]@��t�n_3�`��9jPh<�����V���N��s��74Ab2w��0��9�ƲL�+0S��g��CG��<Ȕ-@�����M8�X|�\@�/4�ޣ'�"�����L@�*�>
z��NeN�W\g��ݳ����$�7��}JP1"�<,jB(q����*<#��(׻�R,��4�t�ӆ�7|��:�1��������`��M��u�-��24I�ɽ�E���rs���pHXn��֠��c��d�ټȰ����e�aZ�u���@�E�s>�а� ��Ӣ�����Q��x�
�pM��EO���#n����*���.wc�Ωnh���<�"�r������0+�}5��J��i�"�W����I��흾Z͕�+�Q����j�ү�;�J�?��,��q��S��K��R�s��☺_����?�~uo�dH��ڵ�d�ɝ��)�bj=3����]�%Y�yMU�1L�4�zi�^��yEZ7��ܳ�7�9�C0U࣊�x'�� |� M��ƒ�����§�b��b9#��r�Ce�'H����[��R���I��z�� ���M
S�Ф)�OGW�&���g��J���?y= �?y�j�1Nʮ}@��[%�Y�6΄kD(>H%Y;?4�c�e�I�7���œ?�g|&�j�������Z#q�+��J�ў_�u�ü�Y>5߫�(6�F�gx� ;녽@�iA-D�{���5l��!�w�����֏�7W�o@nE��\H�q%ϴ���QM��ݮ��í�E�c|NƦ#>e��.��� ����Ш�������� Vl6R�d����槵|&ft�7D�r���قb]�Θ�'��H��>����u_�T�r�'�;���1�=��W�`"ѭG"6���\�,,��ہYBlۮ�l9����T�\�y�C��s�U�y�35��N,��Ӿ��7�>�/f���5MG�mx�/SZ�����忐
�Ӛ��0Իa�����,��ZSI0|8���77�w��x�	J�+7z@�F��J_MA=Au&�V��vQ��T��j��:�3����>+��n���)G���5�y-wI�.�f�;��/��v�m���~Z!� �'�V����Ɲt+���u��FS	��K��GГ�c-�ʡ~�k]_6{�ujUD�LX���	x��OeoI�.�^C�r�'y�s¹B�����O���(�|E����}�7�� ��鄫0�Qr�`6�yb�k6BXO��VD�yOuuCf@�+�|�I�;[>]JJA�Z����P�x���&�e����\��	�U�3�S����_~�\�F����?�6~�L�8m�����XŞ��b��Tڴ�"���g,����G|��N����a3#-���N�����4����?��٭�[�S��P�������w�Oý_�x>��F��"
s����ٛ�k�e![1��?�Z���M

�63#-�M��[�cM��w�(�#����T���I�ݫ���?�,I����O ���[��S��D���vD��uzKQ��T{*�ab���%��aO?�kΓ+|r�?:�y���|�y�L��d=�2Wg2���yo�֝e� �I�RC�7A>�w�Պ��X��ѫ���������m��}��k}��v����'���s�轘���}=3�NA5�"�#�;�S`��#�lUZ���D�ˢ��S�R>T�_�&�Ɵ�@�L/r��mG��=yO� W�KƙZ�t%��uC��@�\2�Z�F��D�/|���G�W�;v1 �w����s�����X@�*e0J�P�_!�Y�!��\,w������ǌ�P�V��WI��Q�1ܕfx�d@'�ֻB�f�cD5�-�}�3^jx�e��$�m�§��5J��^�3_���.�jShL3!2�:֥�eC�ۋz�â�e�0!6��g�;��|�T�ď�/"	���3_<'o�憿?w�+Ɏ�"a6A0Μ��C>�'8���*�א�jHHȈ�|�i���	�s�����[�s�Q���;M_�=;\?.���!�	z<��۞�������R�i���K��BiO����\�Vmi�����s9��;��vcU�Ě:�����eQDsV�?�4[�`��VΨ�8�s�$2���0�uG�/��U�if��q
�S)�����	���ߵn\c�7�է�Q �^Cng��?A~3���_c��t]j�f�{��cH0�ʪ5䙴u����~}�ض^E+<ۈY���6q�����q�!~�6��~��J�)�z��4�=����W������E�UP�!H{��7�y�������ܩ�(��!��%C��f*$��TBw�l�/���˃����yx�8�/��RJɺ�����%� 2��C�
��O�-7�s����w�i$s!�ʖeF�#��m�"�������b��g����k�/�Ҷkd�8ݾ�d�lvD����������瑈��:Z������.�1�n���<'���0Mfkȭ��l���B\F�@c��7��.L��$,� �h�� �`����x&���BU/��K�AA3U�p�?6���qq�b�v2^��k���`}x�h@'��v�Wz#ܟ��p>�Ur�#�<�	��~	B-8>�a���q>f��+e��\fR�쀝��!��5�-x�v�J�x��߂T�
�|��U,?�ΒҎ�1��&�Ň$W]N��2�������V�k;�yu�=�x�=0��7����+��Չ/�o+��E?��Dy�9���6ٻ�����+1���{?�7�̏<j�~"��eV�ه
A&�`��ɳ��.��b�0���:����'Vz�\dA��:���E�X�b	�e�Pbųr�^��'�)���ʯ�b��jւk�IN{�l��վ�T#W(Z�Y�V���eO� ��MW_5��W]�=�	�����z�E��6��Y�M(��Q�H$��1�tv	F��b���$��B��*I,���u+8�rLB���t>��)P�2pP97f{�|��ǹ�����C���}��������YE��*2PӘ��l�7��o�(G��o����&��1��]k�1��� ��A��U���8">��ъ��P�֖�ڐh>{3�g����Dקn�=�-,P�v�#��3�\	2bGk._�u����/�ɏ-$����ٶÛ&~��A�%kk������z_:������GK9����aS���2^�*<shЮKؚ+��{[���1���ʀ�?���4D^�*�욊TE'?�up����+M�s�$�z�ž|�ݩ��e�3�8y�,�"�qh�J�2��/)��d�1R���6���J#�L@rٮ9Wv�5��S�fh̏Qe��P����q�l����b�J2��kQB����[�$~� >~ȓ�&����"������~{�)��%þ����8���� ���`�Ѭ���d��b�C�D��VX@w����.�2kL��k��Ռ()Fd�Y}D۝au^K�n��m�ڼ�Nי���s۷�- a�u��R���8@�r���sA��MK���=���/=�j�@����S��!�����L��,�����IÜܿl��h���
�Cs>o��3�Z����P~*�S��.�R1�>vs7l�t8o��vB-��5�V�:���&�Q�V�R�='7!��Tv����gq�qq�}�T�R��[�6������B���ɤ*���M��.�1�>�sX#�Zj]�ՙ�؏vv����ӣ6N]�뻋����� ��Q���I���6�/���G�Kl�05�H_gT��^s��D.Z����lz��zUW����\D�p����e/�^���F�&^�����!���V)7�q�(�i^?�]��.ȝ��l��-�!�2���L��0ITgd'RٳC�m�������\V���1O�F��L�)��ᛷם;�zϿ�`�<1'��m��*J���K����dc(��Ǆ-�����G� `�cC#�����K4�L�E_k�_'x�I �R�L�|kr��dSt����i˙�&���c��^S��Cр�V�O���r����񁇭��;6�j~�.Z���:OY�W�o��9�h��lBRO�^�5-��!9�DWɧ������*��J���9���&b}HĈ=�#O���!�H�M��!�Ы7�J|ɑu��0K2�/㾤6ᘭ_)��l�=�,�7̴�r����FR��5�j�Q�f4<�
:q��d�j��\�C�A�o��6�Io���ן�u�/}5��6#�KO��%l0 ����bJ�0�2fX�A��B��kl�P�I�/��)�a�K�db��� �����v��u���r�p��=%l����,?�������8��M5&A�/>ڌ	�r9u��߶lm5��2�Z�)
�Ռ����ՆE"���Dgbm>*��I�����*�"i�C��6u��%�)��.j���ġ�Lc;w/
��E[l�j#;��.�?�SU����m�[�c'�]GM�����azw�W��cN�9ǜ��e!^`�G����U�nX�|ވ}�}��,���.g~��	����^, e����TA��=�D.��i����(@����jI���DP�VzTu�{$϶1p<m�<	���U2�L�e��^i�m<2����Y�e]��3��}��TC��7�+Rg�l�R�'ȵ�g�t�'U\H�(-�"R��'��j�P�XE��Ꭻ'���tDk�^kun�@l��?(�	3E{O���� '�v�t����vź����!���aͯ�z*�Vs��P,Q,l`زg�� �M3�m1��z�l�����{f���vih�O�|�%��WΖ�Qk��\<}G �r����9uO�m}dC�������8y4���_T.��x�[>m@E��#�WC�-��=l�m.
L������b�`#<�3P�޸
�;�p���uX�:��чc�ġhr�� ����lf[]�Y���Y;h�X3e)�ٙ�a��a��c3���]ݰV-zf�r�&��S���;�ܳ�����5	 �0�-Eb�w�ߌ����!����='/˩��Ji���8-��& ��
S�w�Bj�
��������[ݳ��!Vfn_��E�oFl�)�\Q����g�i�Y=��������N|�s���TL�TUe��s�᮷��j�5��X5�A�)d�k�FilU����țK��^��1j���M�)��X����^T	F�j6uG��ak��*��^��o<��5���$m���ȋO�/��	<6�MZ�;����6�h��ׂ��_�x�L'���9҆Y��^��3H@� A���͊`ƺy�M��rQ��Ox����^�O���%�=,��O�e5�%^o�=6ݻ����P��p^���!aLY��Ϯ��'��*�
yN7c	�H��!'��z?^�`�.Y����Z�@���Wm���k��8��?�56c����1���6�n&�*dW�`��c������W�^|$�|/�?<&�A*0�N����?7a�������PV���"�r��՜y����ruh�3!/��3f>�-BN���!��/+�f�V����k���l|/)%����	�U�%�x��ފ��k<�M�/_�I�9"���IvS��J���%�s�1`������0�W(�����oJ^\ ei�9��7��E�.%���]~N�ɦp��F��>y���X�R���c�6�O����-{W��[�jt�H���-�o��1�\���_��r��p�g��j~'v�b����X�?��7�@dĺɺ��u���b�z����ଓ&�$C�h�����}o �*Aj/;����!_S�ß���y��+.���&� ��s81
һ9�<�� �[��0���J��D{KtkW�1��q�~{�ל��c��]":�>b���ʦ�ᩏFEwo�͹����4е�2��]�`�a�.������v;���͚���d>��B�H��яJ;��V�Lt�-07������Y�,�����h�����,ŀ�M�����񢨢�Ѥ�1�|(�钎A��K��-���-΃�.os�`s���ߔ�/�@3l�3
�dn,��g���̘�F��wo��dC)���a�s�ȥ�K����i��p��~���w#\�4Yk<f*��	���}d���cl�:��W@�t�]�;x���jX�Edj���^��K�����6�<�Բ6bh�o�5�}X>}�L�����Հ��)[78c*,��	��������+���W�Ią|!62ˑc��伴���xR1M��IK+[j�����Õ� H��p2l��	��5ܱ��|L��߼�SIs�VTY�I���½$Й%���ᦢ���Ě�wpk�-T^�(W��«�bח��e�k~K��o]l�����H�W!`΃��h�*M��7>�}|~��DF��ڪ]J�_��v+1�N�ǯ!���[b��g���˓���_�e���B�%�0�i�ÔӼ{�j_e3
r�=t�����M�
�Q��*��"��l�F�$޳ʆ���V�Z88�(1���GK?w�k��f�R>�a�jc�j�f�@+1�9�<3����hZa��Z��>gcͬ���f#R�!K�M��@�,�֫ �ۜ& ����g��I�CK�`q3f'�e(�H�V�H�K���.>��`�+!�_O}�@}�y�YxS����L.zD���a\dl̋���
��^Y���)�_+���Ꮀ������ﰑB$��ځ9��s��>6,�*�x���)���j!�	�	`.��4՘�}�/9�0+~Q1hu�����������Ou�X >dZcP7#MI���>r�'�F��A4Ć�(��]�r$�l��5~���a鼢]�@	.��h�z�6k���V:�K���ԉ������<a�,��J(����I�}0�f���*2u$�����N6�j��h���ן��h�+H�C��I'�1�_czs�#����FS�x�v��
g��d ��Y�D��C�08�������2#��[��I��O�|	l�g�O�V�.�8^0ag�ͅBl�A�9�'��F�e��L���I~A���!���p(���J`@��gT\PN�n���!Et���I)���.����-��6!܁P	��~������@�8-�*�[���[ƽ W���2��V�twdF��ΫT3��^���x�r:�1�A���x�w�S��s��^٤C���	d��z�Pv܆�I�͍������h�1��]�@p�nv�"O�S�k,��d����ҵ9|3��Ӈ���FX#�g� �29���iCQ�哥���?e6v�CaHwjǳG�X��G�o�/��i��k5��ͽ�N�ȘWX�-ƪ�R���Yi �_3cR]{\��p���y�US	[�w�!~��|$��Kgd5߸[�-��@�yG���i8����#;_��������{d������8�ݢz��۾�@��];=�������y��:���gR����eȀ8��dI�$C[��W�ѻk������橡M\���l��t��a� g�r}�d��w�$?�	~3@��om��2�{����kP��K�r@��Ԝ!����y��Q|��`��9$�ؘ��f�Sz��:n{N��l�F�_��Me�;�J��}qt�'"|�_u��LE0Yn��̱ho�5#gG���~�*5<��%e+�+1�P�A�ov��[�ng�8d 8�"q�;Ǒ��m�y����Q��^�:�r=�4i':�z��0z�Gl�E�G�\��_y��Ry;�~��Dm�3M.�إc�X���j�V����Fx�Ϳ�T�����dki�_4ο���=W���Dn�C/	6N>n�'��G[X@M��?u�2Ł|��)��v��̨v"zǏd����z&�pP=x��}ґ��E4�̽E>n1��$|��mDI.�!c���=��6Z��'�}�ӸH�hB�,�����y�܋Ow簀rsp���Rⴭ�������Fzž�A���f]�P�i���f|>���E۔�i��+��'5�2bz�5�ص��P�m�Gt��G"��6��.����c�h�:#�E�YV]Z
�� R�,-�S�·A%E�65�!1���O����R�z�c�ٍ�m��n�S�(���eO��b /M��c?9���km�h.�7���;���gmu��+_·�f�������dj*:m'6�Ks������~Z��}���j����+v�����<#�-����橃�es�ت��t�n�q�B,a��YB�]�n�ݯ�T��|��*�Y9�-7��}�}�}�@�1j�o';��j!fr۩�$�cuN��.ww0<���*Н�[�{�<����I� �JZ�W���kF�w,�4��X�����4��h�k��a,�O��.s �Zxdk��X,˨�N�����GCl��Ƽ	�~�~��;���i�b�ά6��~�;^Б���"�nu��������-g��K@姎<���|�Zٺl��6�dr��K߮$�m3������L��.]��"�3��<4��iҬ��nJT��8P���y�ݝ�\���!ktŒ�`Z.�7V̚ƃ3�D�e�������5���M�[2�)t���X���J�x�OO/��,����C���'��P}x9��7:��i�c��x_8� �^+�{���[w�.s�y����a��>�[�w�Q�xй�f�ߊą���Csz�L�ziw�$7!��Ъ�
�O8�dR�Ӏd��sHH~|�:w��.hKS�����+���z$"8������0�}O՟�Qq.�x�9���
k��y1--A������}s�I�"�D�OT�J4.�HY��g�I���V7꽪>R���ݎF0��~�ꅖ���4M���N<u3���>��^`& k���:!�ꡭݠ�5��^^�jU�-y����)>�	�<�i��q��{�qj�<cK������9��J�ؕklѺz]��կ������[�T�)C��*��B��M{��5#,�>�Ξ��T-�(��GU]l'˖qM�|���O�8��b9�np�k�h��l�I���yO}�O�_�~�U���\�����PD�{߂�g!��ۍC)onu���K���x�qu[���9���"m�0v�366D�U�b�?!�=�!��'F�_�q}t�	�
_�O�N7,5�
X���VYj�:ۙ�GrN3+��*[�Ō2�m�SҮQ���/���V� ~�V��\]BC!v�B&�b������Z�C3z?rw�
�˂�o�og�!���n�N�T���������G��T������2��tW��xe�焀Ah�a:FEΈg,W�7��x�j���z 7�0|+��Ceٞ2G�J5�X�wK���*4c�z���S�EW۬#�+D"L����*�P$qz��3�G��-��ɒ$���ԇ��u1̑�%q}0�Dc%/�7�~QOf�$&����E2WD���/EӰ ��jcS�3����&=F<�[�,����^��5,�Y��㩴�+����q֍����J�������/�����ȧ�;��I���V��v�"}��'r�:[m�5���`I�yi���l�oKt�O�2 Ȅ�.���V�K3Y;tW�ST!0�a��#�8W�b�����"�!-���k�Ρl��	��c�snw~�]�n+�eh��.�;��6�7�j�U��G��g���4i�#3��GA�G���&���׸��\9� �R��E�5�b�A���Py���}�R��A!�y�x��<��e!��n����0�WtX���{���x��)��Y}Sj���l.����8���vB�@��_�PM-<-_r�j@f��1U Wc�ǌo�~��j���]딕MLw�='��s&���Fm{�#]Um���������f3���I����F��٬�7J��ر�-�u�7S��(ef�RmÓkO��mI�/~�!hc�0���Y�m���Y���і�=o�;	��p�"�{�])eՋ�KD��Fڱ$��O�CpӞhv�	����Iޝ��^HA?��z���3+�wА|�̏��]��u[�P&�%Y�{&����MR��s�q���ã�g�K�8`\��A�t�TW���z�V����&�����x_W���ٕV�w�e�&���"�xӥ}?�t"�HCV�ȋe�� f��;�໥D�lx��B���s���Y>�PZ�����]��^�VV��~	LT�����`��(��B�q�?4f�h�N�D�)�NXc��¹�?��Ƨ�����h쥔�u=����@�l�~V3�d�=*�P�@�](�kȨ�Yl�>�1m�/^�[���.J�^m!U7���c���]͢0�T��0Xr�0!�
 �~*�*E`���c��[��zF�+R/`���eX R7�E�6b~wrB�8��W�?�T����?�O��r����!]L6V�<uy�l�4����[�]%C(UP��E7�+�pF����������e����F.�%E��~[cQ���a�,��|�dz)]���7f,lr/STN$�_=��,kpR"�6�(�
�����!��7:�%�����S;�U�	��>,>�a��9���ڡ��⌍4g1�����6��������1L���
��Iцt"��<�~;�%l���f`^���dby�3�6� �NF�?W��=�����/I�,+�C��h����H]����=V'7=�����<8��y �=���ؓ3���ID�O�����5�n�g��z+�?����#e��U��f;����r���#��a���hKNou�Վ�2�����(�jq�?���@Gs���կ�6��uM��^�����4����k�3&X@hN��OkD��[AOK�/7�n��܎~��^۬�9�?yӅ�r�� �@��Ȑ#�W������nR����GX��� A��r5�8�Fi����鱨����fXS�G�ӕwGj�&ڱi}�|��Ar��#����x}�����9R�����&<�T=��������� ��p�f��f�m�f �����Ub�]�,�y�a]-�^Z]뒷�<c}��-�q�P��w�f��#�Xu.���,B�XPRM��j=�3H�MZ n>����]����I���U���[��C�qЯ�)�MaP7E4����*�4�y���r|�H%��L{�F�Yj=7���&� ��1�Q��ʱ�br���ë��հ�UĆ4ۤ�wb��CC^���l���ȮV�j*D���q|�%��ŋc���L>E	n�%�C+ͻ?|e}8��Phl���U�N+z���nٽs�D�o�?->� ��N*�{����]	�Z���EF��t�g� ���f�Ӝڗ�'0m|$����P�����+(l������b����z��@r��no��<���Ms砀�Ο&�t��)\����ӽd�0j���*FLNC��H�+C~��>�V�7NUҰF'�R�mo���I��|:To���]�j�z{�<��k0����~}�@�fq���0��P�߼ja�=2v��"��ao�M腆)�6$tYW>��v~e��*Q�͇�@b�<I*�ԙ��z�4q�yV _�쑗��h{�ͫ����ϱ�0��$���UՓ��l��Z���B.��2��t��Oo���^�D�Y�ۿu�?Po�(UG���|먪\Jf1}*�ɖ3&��!�����Ț�����m�	1J���[��U�0;���(K]��o��z�xӝX�lҩ_/f��
�<t�8ɼ� ������4:7�pK����q��YD)�+��v���H�g��ָ�����y7f[����%:=|��%;�x��[�b�
5��,�^��ݻ�A&����Y�'ՅV�I���Ϟd�U���z�}TY}����;~\�����,��:�E����ܻ�s2�$����+.1_��6�D��݃����1G7�t���<I��� �o�}0�׼�@N�@�l�����x��m��%p6#׷�4Y���*��rc��Ж����E0�@?�M�a���@�p ��Ӱ���+QcZ8��;�W��t~���E�1T�hD��+:3����1�Ϩ��/sj�qTd�s�u	���
Q\u����!b�\?�'�����x~�Q�\�%�l�XVzy�A{yd���-i�`�W�3��+H-����2_P�j�U�d	t<t�}^.��=R����b����ȍ�vԛ�.qq!�L��?]w�eu0*f�oQ�a������&��C���ic��&�]2ԛ���h���$Ї�a��S>ˈ74�eu����+�qk�^�]�s���9��|��ނ"��#�5N_����q�2^=�H,ȵ���Ԩ]��D&qV0u�wg�;��Л����Dŀ�����]��rC�M��u�8�N��yu�B�I�9���Ma��N��8HZ	�}ߏJB�Q��0�x[(P�z�3�3�J�-���"��DObD֌R�0�S.d�vĄǲ��Gt!!�/L|2���\���9���:��o���G���|6'�}�EE~Xy�wA+h��,s|�i�$#���"4Q/Q��|3�}�;{�Q��o���+���oc#5Y��?�7�:@ۘ��j!1��n�2K��-��(���#�8�9�� K�9䘁'���Sw�Ȯ>�}��o�: �hҋ��Bf��~�-��MJ�C�Dd�������.�:�r"s!%�)���g�*��v��P����7����� ɑ1º*�T���ƃ:�X��}��1�JO�I5k^S��DD��1�ل]�+*^�z��>j���H: I{�5�w�0�ϱ����ʥ�m��3����j��Ɨ}}�����h�Ze�h���IF$c��۝x�i��&"��`S��'#�C��{��Tٽ;����p�X��:V����H[l��E�����g��K�j�j�YXjX�C��DK�ʈ����H���2��C��B�To"^��Y�ކY�[�dV�L1��|e�,?�E$s/��<\��X.���dLqzK�|~�ش�ϴ���x�W�pp��ܝ�)�l�=_��̬�ǋ� ��֠	-������_*q���2����b94^�.�統��g���s�ǜAzaһ�s�����ڑ)�Ƣ]�8?�<�f�#�`�TS������paj/��N�@kY���}�8}�,�R��K�"�!	@�fQ�ӯU�P[H_"_�-�{R^�&��-@w��d��bo�F��Mߵw:��v�R��!��l�E`�F0��	��JG)H|�Z�^@�oftS�j'�ؖ����ߋ�x��X��iW�#x��a�6H �-�<�7l�jD镥e�2�w~,���Gw�]�`���.�0���ɾ?_Y�w/>�Ԯ�5���{���(=�CD����1~��}��X������S-e����Gהц�����1݁��5m�a�0�}�W.��}/e�0F��|�ܣ7���QL��z�7"?6.��s�S���*�5		΋߳��Y���8�ί��+��Y��?q��G;a�V�|�[ٽ3Hs&�ʐ�47�ݗ��<�Q`�˟Q��)��J���+f��1���e�NȳV7�i����$�hܟ�g�N��a����_]UȎi"���y]^�$~roW��)����EȮ�u;���P���M����L
�$�0��R���I_���>>�K����I��{�4-�Nv��;V������nPB.��v� ����a ���*�9&��-&1� �b�����_p���I�1l<�
:�]�qmp���q�q,���?{��
Rz	�c��L�#�m����G�<��h.�3�^'����^�gk��c���["��n���i�Uw��vW�W]n���ކ�:/�i�&jp��+b[�7T2�[���#����Y��@8�u1p���ZW�̉|G����8�n�
�3���a�������q�x3���� �wb(n�
E����0n�~7�W
9������"!��/�%P6�Kj"��o��FB0u��H;TQNy�L����6��`��� fw�H��b/	�I�Wc�$��}��*M�	Gy��[�+�;�6q��{>�CŘ�߷��8��>�P�]Y��m�K�@4J��4�q"U��E��3�\�+��ߐ/q��H-q�R �mM���S=6z��I���y-~�;O@�^�ε�PO�������"\6Ef.3��|�uis?0c���	��EnI��in䙭~\��K�PQ�TZBQ��/܌0���~o��1i��tfS��DP k�-�	0�r��/�f2�.S��]iA�\�( +�D\=�ڃ�C&K5�(��>t�v������RX1��x������p�pպz����8��ʄ����N:�*<�K�
�
���J}NįyZ�3eA�!�����)p鵂���[O��&L��MD�u����:����@�7��|8�_�������WcY�R�~�y������t|D��/���l��F�f, %��ח��=���B��+ojw	a�b_4+�	��� Ɓ/PiX810���Т�/��5`;H 4�C��k�1��&�����;�=��u��T/_�U��b�w�Q����#������xr��:f��� ��sISr�g��:�^;��Q�1%5��aΨ�����Ӻ���߹Z���="i��7_��a�*]���r(`���g�U��ep;k�����c���l�J�N�-Y/���ߟ�5��tXf\��u�ѭs f*��X��x>�Ii���?�/Z�˼�"�hϕ����\�a��з��(4	L�u��o6�LY㛊*�2�"&`��V�ғ�X O^�8��X�;�t�ˊ�Z��S,�O遮S�Ch�^[P���z����Λ^08��x#H���([@��h�gp��i�e'�����O�l�;^Q2���~r�����G�V:���9�Ҥ�Y)�m�P�����S�����§���:�V��:mQ)wץz��x���x0���8��/oQ��k�V#�ѝFPG���d�����Blq��,V�1�9��$X��P�ia�4����<P�{�a��G�t��'����E�1,���]��]�\%0�|�?�Ѳ܈=��t_�,��Ή)0�A5FS�ۘ&�:'��l�&�ѻ�����$��8���y$_�i)�����|*_Xu2�7zMT��F}���eY}�w.L;�/@�w�G�E�p�f�J;�Zۊ�"�^��Xf��n�سS������M�;r+H�,��҄�8�:+��$�q���Y���e߽���
E`S��0��C}/��+�K�h���"��~W���:�Yi�Dv
��������\�Yp��0-E�)�o�/�>�O��;F�6���/�t4�`4�,q��!�ZT��B���WF��!+���������پ�8����"�dt�����	R�U� �P�8�>ڮT}��%%u����|�eq��՘#RGE!:�"HܚD�v�~x�����z~��J�o�>K�Q���Eb�%��c�Z��
�y�N�i�.Y���x��57�@��F�j�WER����}Fص�b+�I�^h��B���W׿E�^�4Q���"�8^�`�݁)�g�E���B0c������z�I6�|A�oU ���`�4w2n-O�w�X�z,��0ҊVjN�	_-.R>@-�ź~E��1ӄ�P%|y-���Zӎ�u��S.]57&Z����ŕc�0OB� J��E�}�d=�ϥ�Mr:$kO�)f�f���w���0q�/H!����Yʛ���Y��U�ƌ��AG��η x��lH:2��l��]��C/���j�6�rw���Bio�B"���1ʊ@�P�~_�w,\�ʱv̉%a�5]����1�p�.��,$�=)!m_ܯ0E�l������8��'kdU�Q�|��i�Vۙ5���M�*<o[��}zш ���xś㔴ݪ�sjv?�ί�UG��%����q��P�:����Ԕ�)�8���I��dn�.���ݫ+<�3��D�Ix\¤\�8b�ȶT} ��5�̻s��D�G�k�O���P��n�CZ��,��MD��|T-�p���O��L=a�T�d��Y�
/��}�gS�<����lBX,5��������E��p�8�k<�����2��1̘��^Î��HG,��i�w�7f��I�p�e�N^��s�	�{�|�H�hr0��D�m�]u�=d�x�ǵ����ǹ���(�hȧ}���0�����+YmW5�7�����eC���	qS
[�%츾�^�� w+\�i|0ԙy���/��Ox����~�$��A�L�rzU$O���'	�5��D�����t�=J4b�Ԩ��,~��9.���U�8�����;�h'>� ��!d��(�h����9J^�yf��~��������	�1|9���u�q���b�i�[{��{���U��k�E��H�$%���(��q�l�����@��J���_y@����vY�T7�U�>G��3�|��-Ϭ�6?��%��iL*���#g�X������a:ڭ��I�e��o�%��8ډO�-(��;�k��=.q'e���F�2{1-)N谳7�xbiFC��̡���j��ą��a������a�qމ���@� "�"-�`�6Y��Ƃx���6$Ղ�y�]�%�+��y-5 �0O�Qͯ`z�yFf5r�z�m��{�V���ښ��\�f�u���2��7�A���b�X�_�����F�@�u�:���䐿J��VD+��>	8UM��V�c��"Z���Z��&9��:�C�PK   �e�XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   mk�X����  �?     jsons/user_defined.json�Z�n�F�A�� j��ys�Ib c���b�u��T(i.	��[�d�6/����M7O�u�������2N_L7�X�bʋ����X���g��6�^������7����ޓ*l򢜼=���ޮ������r_��,�U�X�j�n�:��y��bg�~�R���!%F�c�,�i����s���4�|�/�['��_��N��E@�+�x iR*��9ުlY���ү�F��gxa?V/6E	�X��Y���ߧ���4_-�˼\�j_M&`�����Ss�lo��Ҧ�݀G�Y�\W9������v�U��+�	<#��G�:)����[�/���fa]�W�={��t�Ǭ��ay7�n�op�.޼����a�(�7q׽��+G���]���6��*�1ES������e�6��Ӡ�J�(�+���۠t�	��4m�<�$��ߦ�'��M*:.�OX?h�Rt\��~�6���?��m>�g���؏��(<�����Sd��P$mZ:w���M,�������js���D�EK���'-�(Zr,l~�EK��5��5K�D���m�5Y{��Gms������M���A��2��n����	�v.>��^��t�����b�K�D�'�(^j$*p�]�������
��?�.h���Lr�(�ZpęN�1�ww�Z�ci�`/�r�u��;���:
=�VC\/�Zv�ŦQ�%�u����w����E1/����Z�*_�no�U��M�o�@���g��d�zS�0�cz+��4졇[�"�=E`����c	:i+^���go��ؼ����\M���uAu_[�.?PT*�Hr
CVX�	�����Fŕ���WX/��q �@����� w/|%Br�-'��$��"�B�&ce�w%j���2�I��ʰa[���ΈT�̈�`x�6D:F݁75��Mb�7}�{���(�Tm�����p��B����擷�ueWe���e,Ve��[g�r����!�F(�WH��!��U�Yc�-㌤VGD��L	`I)�B���I�8�&*S�+�E�Q`�9�%��A+Mf�4F(?0���Ϗ ���!�^������GL+��{��s&����.�[����>�����F<�/_�#"�4�/����M�4�ޗe4�@ŀ��F
�r��8B�`Xk���s�}.����S`��N��L'gt��No������0(YX��m�� (A����Ѳ�G�{����(�q�l��!*�G<q��Ω \v@b/q���}����A;�4q�(�4i� ����榁�!��$�.����)�s�iM��A)���0gW�p���S�>�]��X0#Mۅ��=�@=��M޵Yr��KX0yU��j���"_�[}��1���6��TrDm�ZA�q� �"q�f�[���Lk��J/45��>$̈́���v19����֯�f���քΘɤƪv2�w�z͈huW��v8h��@9��Î��9� 8��^]��<0S�v�0�IL��g�j�;�R���df�abЏ����2��������_u�����nw$'�T�|rȝ����4��ݖ�L
�m��83|Wv	��h��Ȇ�4�%�9�̾z�S�F!�e@<���fA~L\(�SdO�(N���~|:w��b@FX�tuc-�^��B������$xd�1�@P(8`��5�yk�x�t���G�x��`fT+pVu��)"��@.G&|x��ߨ�C��]4D���OQ-��z����?%C�g)�;JV��M�Bxh>��HÛA	�-����t�?آ��I�M�˰Y�Q���Ku[�$AA+�ht$;+�\PV����K��A!�l�� M������-���N�QJA!.)��лE��ܸ����hQBL�U�Ǐ��2��$2#���γ�l2pXc��:ԐC=t:��74��U�����|�ڲ�ւd,cB6�`�-�.��͎#78����ԛ4�7� 6gD����M��q�Cr��z�55�1�š��3z���3�1A�9�D������Q&�O,t��o?���Y��sWw��(#��c��gd t�Ѽ��@>��5�2r5�s�)�;&t��C�;���|�����ǜܺc�`"2,�,��5`]'#�6(�NP�j��6�)JWݧ�ʞW�U�Eo2f�h���ԦB ]@EVi�T��:kn]�O:~�V�h�C�@���
�|���@�/&��V���J��D�Sh<��ۄ���Sh�ퟮ����,�^�l�-Y�)�P|%�3I2j���r�n�c�(�?��E8���?����c���>_C�=�o�
`H3r���"��q�g͐$�ZΔ�8��B�����P��A�<��D��$y�T
�ߓ^7A�{�[��/[��	�ߐ����W~�|�`!���/�u9�!_}O��j�[�nݹ��T{>(o�Ϧi�/�7Y�������ۍhn���޴����U�)p������]�3 /���{(r$T��-�匏�*���2�-�q?�#�r2����OC��Ә�I�(&�iB��
i�t��'�Nc;*�L^W���^�cϚ�	2 �Tm4ȼ��PG�$$�e8(I�X�?T%��P�hО�@l��i�B�)�u�l�v��Q��"��i}���ա��9D���X�!O��z=9�w�x_3�ia�������jWu�ڝg��9��&PsΟr<E0��Χ"	PU%ED�k���E�CS��Q>����;�s�_�;�uĳ�x���:���PK
   mk�X1}��J=  b                  cirkitFile.jsonPK
   �h�XWC��)�  � /             w=  images/093f54e3-331f-4155-80d0-fca9fbcaa25c.pngPK
   bi�X��/F��  ��  /             � images/24a65fc6-6c28-4ce3-80af-2bdea9058a0a.pngPK
   ;j�X����7  �  /             � images/2b66d102-ef9e-4dde-8ee7-817842500f7b.pngPK
   �f�X�zm�B	 �
 /             r images/4b3ada2b-268c-4f4b-9789-7d2b3b5aac60.jpgPK
   �e�X����+  J  /              images/5644ca41-1cf6-484a-bb07-c2f9a6f5b19b.pngPK
   �h�X��_8
  3
  /             y- images/57489f55-55cc-4ea4-8258-f1cf3d9c722d.pngPK
   �i�X�z��kW S� /             �7 images/65d233e5-7445-4b75-a6a5-2d8c2ad1af28.pngPK
   �e�X����H   C   /             �� images/8e6e9996-4250-48fd-a42c-980e5b13088a.pngPK
   �e�Xi�={L  V  /             K� images/938ff297-106d-4ecd-b830-d3af457c8fe3.pngPK
   ;j�X�&�}[  y`  /             �� images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.pngPK
   �e�X��) oj /             �* images/9b962a8e-14b5-4317-8666-1954827ef6fe.pngPK
   �e�X�/ w� /             T images/b50388db-476c-4829-8b73-5cdf8357e0ac.pngPK
   �e�X$7h�!  �!  /             �a images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   �l�X���k�� �� /             Ń images/c6c89cf8-e908-43a9-a5fd-b5d85c65d9c6.pngPK
   bi�X�ة� � /             �D images/ca60ea1b-712d-4ba5-bcf0-f1dd45701dbf.pngPK
   �e�X~��a� ٮ /             �^ images/dc707dc6-8489-41bb-a5bc-77a0670f90d6.pngPK
   �i�X�|�	  	  /             m images/e1d4e862-170d-4bac-8b1a-e4319ef50e6b.pngPK
   �l�XS�X'  S'  /             � images/eb6b75ee-ffd7-462d-b06c-ecf58549be32.pngPK
   �f�XK�h�� 6
 /             }D images/f2a2d8b8-8493-40f2-a2f8-368c45be6cc3.jpgPK
   �e�XP��/�  ǽ  /             �M images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   mk�X����  �?               �� jsons/user_defined.jsonPK      �  #   